************************************************************************
* auCdl Netlist:
*
* Library Name: SMIC_MEMORY
* Top Cell Name: S013LLLPSP_X256Y8D8
* Version:  v0p2
* View Name:     schematic
* Netlisted on:  Thu Sep 19 15:16:10 ICT 2024
************************************************************************
*.BIPOLAR
*.RESI = 2000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH Tie_high VDDP VSS
MN18 net15 net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 Tie_high net15 VDDP VDDP P15LL W=4u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL TieL VDDP VSS
MN18 TieL net15 VSS VSS N15LL W=4u L=130.00n m=1
MP18 net15 net15 VDDP VDDP P15LL W=2u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_inv
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_inv A VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
MM0 Y A VSS VSS N15LL W=nw L=nl m=1
MM1 Y A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB BL BLX DBA DBAX DIN DINX VDDP VSS YS
XI7 YS VDDP VSS net81 / S013LLLPSP_X256Y8D8_inv pl=130n pw=800n nl=130n nw=800n
XI4 net81 VDDP VSS SL / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.2u nl=130.00n nw=800.0n
MN0 BL DINX net58 VSS N15LL W=2.8u L=130.00n m=1
MN2 BLX DIN net58 VSS N15LL W=2.8u L=130.00n m=1
MN3 net58 SL VSS VSS N15LL W=2.8u L=130.00n m=1
MP0 BL SL VDDP VDDP P15LL W=1u L=130.00n m=1
MP1 BLX SL VDDP VDDP P15LL W=1u L=130.00n m=1
MP2 BL SL BLX VDDP P15LL W=1u L=130.00n m=1
MP3 DBA net81 BL VDDP P15LL W=1.2u L=130.00n m=1
MP4 DBAX net81 BLX VDDP P15LL W=1.2u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUX8
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUX8 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6]
+BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] DB DBX DIN DINX
+VDDP VSS YS[7] YS[6] YS[5] YS[4] YS[3] YS[2] YS[1] YS[0]
XI11 BL[4] BLX[4] DB DBX DIN DINX VDDP VSS YS[4] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI12 BL[5] BLX[5] DB DBX DIN DINX VDDP VSS YS[5] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI13 BL[6] BLX[6] DB DBX DIN DINX VDDP VSS YS[6] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI14 BL[7] BLX[7] DB DBX DIN DINX VDDP VSS YS[7] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI3 BL[3] BLX[3] DB DBX DIN DINX VDDP VSS YS[3] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI2 BL[2] BLX[2] DB DBX DIN DINX VDDP VSS YS[2] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI1 BL[1] BLX[1] DB DBX DIN DINX VDDP VSS YS[1] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
XI0 BL[0] BLX[0] DB DBX DIN DINX VDDP VSS YS[0] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUXB
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_nand2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_nand2 A B VDDP VSS Y pw=1u pl=180.0n nw=1u nl=180.0n
MM3 Y A net26 VSS N15LL W=nw L=nl m=1
MM0 net26 B VSS VSS N15LL W=nw L=nl m=1
MM2 Y B VDDP VDDP P15LL W=pw L=pl m=1
MM1 Y A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_SA8
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_SA8 DB DBX DOUT VDDP VSS ck1 ck4
MN4 net85 ck3 net94 VSS N15LL W=2u L=130.00n m=1
MN0 DX D net85 VSS N15LL W=6u L=200.0n m=1
MN1 D DX net85 VSS N15LL W=6u L=200.0n m=1
MN3 net94 ck6 VSS VSS N15LL W=2u L=130.00n m=1
MP0 DBX ck6 VDDP VDDP P15LL W=1u L=130.00n m=1
MP1 DB ck6 VDDP VDDP P15LL W=1u L=130.00n m=1
MP2 DB ck6 DBX VDDP P15LL W=1u L=130.00n m=1
MP3 D close DB VDDP P15LL W=2.8u L=130.00n m=1
MP4 DX close DBX VDDP P15LL W=2.8u L=130.00n m=1
MP7 DX D VDDP VDDP P15LL W=1.6u L=200.0n m=1
MP8 D DX VDDP VDDP P15LL W=1.6u L=200.0n m=1
XI53 DX DOUTB VDDP VSS DOUTBB / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI54 DOUTBB D VDDP VSS DOUTB / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI74 ck1 ck4 VDDP VSS net137 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI73 net156 VDDP VSS ck6 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=3.2u nl=130.00n nw=1.6u
XI71 net152 VDDP VSS ck3 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.0u
XI77 DOUTB VDDP VSS DOUT / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=3u nl=130.00n nw=1.5u
XI70 ck1 VDDP VSS net152 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI72 ck4 VDDP VSS net156 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI75 net137 VDDP VSS close / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.0u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_tgate
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_tgate A EN ENX VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
M0 A EN Y VSS N15LL W=nw L=nl m=1
M1 A ENX Y VDDP P15LL W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DATAIN
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DATAIN BWEN CLK CLKX D DATA DX VDDP VSS WE
XI136 WE net122 VDDP VSS net77 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI4 net142 net126 VDDP VSS net82 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=800.0n nl=130.00n nw=1u
XI3 net154 net126 VDDP VSS net87 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=800.0n nl=130.00n nw=1u
XI21 net114 CLKX CLK VDDP VSS BLATCH / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.4u nl=130.00n  nw=1.4u
XI5 net146 CLKX CLK VDDP VSS DLATCH / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.4u nl=130.00n  nw=1.4u
XI39 BWEN VDDP VSS net0206 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI37 net0206 VDDP VSS net0207 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI31 net0100 VDDP VSS net0104 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI35 net0207 VDDP VSS net0120 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI34 DATA VDDP VSS net0100 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI30 net0112 VDDP VSS net0108 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI29 net0104 VDDP VSS net0112 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI28 net0108 VDDP VSS net102 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI322 net130 VDDP VSS net106 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI321 net106 VDDP VSS net110 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI320 net110 VDDP VSS net114 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.4u nl=130.00n nw=1.4u
XI22 net122 VDDP VSS BLATCH / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 BLATCH VDDP VSS net122 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI143 net77 VDDP VSS net126 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=1.0u
XI323 net0146 VDDP VSS net130 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI19 net87 VDDP VSS DX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.44u nl=130.00n nw=720.00n
XI20 net82 VDDP VSS D / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.44u nl=130.00n nw=720.00n
XI15 net154 VDDP VSS net142 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI36 net0120 VDDP VSS net0146 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI27 net162 VDDP VSS net146 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.4u nl=130.00n nw=1.4u
XI9 net154 VDDP VSS DLATCH / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI7 DLATCH VDDP VSS net154 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=1.0u
XI25 net102 VDDP VSS net158 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI26 net158 VDDP VSS net162 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMX8SAWR_BW
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMX8SAWR_BW BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6]
+BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] BWEN CLK CLKX DATA
+DOUT SACK1 SACK4 VDDP VSS WE YX[7] YX[6] YX[5] YX[4]
+YX[3] YX[2] YX[1] YX[0]
XIYMUX4 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6] BLX[5]  BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] DB DBX DIN DINX VDDP VSS net86[7] net86[6]  net86[5] net86[4] net86[3] net86[2] net86[1] net86[0] /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMUX8
XISA DB DBX DOUT VDDP VSS SACK1 SACK4 / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_SA8
MN1 BWEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 DATA VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP1 BWEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 DATA VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
XI14[7] YX[7] VDDP VSS net86[7] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[6] YX[6] VDDP VSS net86[6] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[5] YX[5] VDDP VSS net86[5] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[4] YX[4] VDDP VSS net86[4] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[3] YX[3] VDDP VSS net86[3] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[2] YX[2] VDDP VSS net86[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[1] YX[1] VDDP VSS net86[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[0] YX[0] VDDP VSS net86[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XIDATAIN BWEN CLK CLKX DIN DATA DINX VDDP VSS WE / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DATAIN
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_BITCELL
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_BITCELL B BX VDDC VSS WL1
MM2 BX WL1 BCN VSS NPG W=150.000n L=175.00n m=1
MM3 B WL1 BC VSS NPG W=150.000n L=175.00n m=1
MM0 BCN BC VSS VSS NPD W=220.00n L=130.00n m=1
MM1 BC BCN VSS VSS NPD W=220.00n L=130.00n m=1
MM5 BCN BC VDDC VDDC PL W=160.000n L=150.00n m=1
MM6 BC BCN VDDC VDDC PL W=160.000n L=150.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcellredundance2x2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcellredundance2x2 B[1] B[0] BX[1] BX[0] RWL[1] RWL[0] VDDC VSS
XIBITCELL_0 B[1] BX[1] VDDC VSS RWL[1] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_1 B[0] BX[0] VDDC VSS RWL[1] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_2 B[1] BX[1] VDDC VSS RWL[0] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_3 B[0] BX[0] VDDC VSS RWL[0] S013LLLPSP_X256Y8D8_BITCELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2 B[1] B[0] BX[1] BX[0] VDDC VSS WL[1] WL[0]
XIBITCELL_0 BX[1] B[1] VDDC VSS WL[1] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_1 BX[0] B[0] VDDC VSS WL[1] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_2 BX[1] B[1] VDDC VSS WL[0] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_3 BX[0] B[0] VDDC VSS WL[0] S013LLLPSP_X256Y8D8_BITCELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192]
+WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182]
+WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172]
+WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162]
+WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152]
+WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142]
+WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132]
+WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122]
+WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112]
+WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102]
+WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92]
+WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82]
+WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72]
+WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0]
XIS013EELPSP_0 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[255] WL[254] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_1 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[253] WL[252] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_2 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[251] WL[250] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_3 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[249] WL[248] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_4 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[247] WL[246] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_5 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[245] WL[244] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_6 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[243] WL[242] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_7 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[241] WL[240] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_8 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[239] WL[238] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_9 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[237] WL[236] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_10 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[235] WL[234] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_11 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[233] WL[232] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_12 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[231] WL[230] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_13 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[229] WL[228] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_14 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[227] WL[226] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_15 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[225] WL[224] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_16 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[223] WL[222] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_17 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[221] WL[220] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_18 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[219] WL[218] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_19 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[217] WL[216] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_20 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[215] WL[214] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_21 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[213] WL[212] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_22 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[211] WL[210] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_23 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[209] WL[208] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_24 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[207] WL[206] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_25 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[205] WL[204] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_26 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[203] WL[202] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_27 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[201] WL[200] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_28 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[199] WL[198] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_29 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[197] WL[196] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_30 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[195] WL[194] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_31 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[193] WL[192] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_32 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[191] WL[190] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_33 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[189] WL[188] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_34 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[187] WL[186] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_35 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[185] WL[184] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_36 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[183] WL[182] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_37 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[181] WL[180] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_38 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[179] WL[178] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_39 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[177] WL[176] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_40 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[175] WL[174] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_41 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[173] WL[172] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_42 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[171] WL[170] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_43 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[169] WL[168] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_44 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[167] WL[166] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_45 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[165] WL[164] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_46 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[163] WL[162] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_47 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[161] WL[160] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_48 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[159] WL[158] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_49 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[157] WL[156] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_50 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[155] WL[154] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_51 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[153] WL[152] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_52 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[151] WL[150] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_53 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[149] WL[148] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_54 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[147] WL[146] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_55 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[145] WL[144] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_56 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[143] WL[142] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_57 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[141] WL[140] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_58 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[139] WL[138] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_59 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[137] WL[136] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_60 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[135] WL[134] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_61 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[133] WL[132] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_62 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[131] WL[130] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_63 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[129] WL[128] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_64 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[127] WL[126] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_65 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[125] WL[124] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_66 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[123] WL[122] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_67 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[121] WL[120] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_68 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[119] WL[118] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_69 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[117] WL[116] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_70 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[115] WL[114] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_71 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[113] WL[112] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_72 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[111] WL[110] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_73 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[109] WL[108] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_74 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[107] WL[106] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_75 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[105] WL[104] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_76 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[103] WL[102] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_77 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[101] WL[100] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_78 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[99] WL[98] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_79 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[97] WL[96] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_80 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[95] WL[94] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_81 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[93] WL[92] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_82 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[91] WL[90] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_83 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[89] WL[88] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_84 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[87] WL[86] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_85 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[85] WL[84] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_86 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[83] WL[82] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_87 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[81] WL[80] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_88 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[79] WL[78] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_89 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[77] WL[76] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_90 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[75] WL[74] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_91 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[73] WL[72] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_92 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[71] WL[70] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_93 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[69] WL[68] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_94 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[67] WL[66] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_95 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[65] WL[64] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_96 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[63] WL[62] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_97 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[61] WL[60] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_98 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[59] WL[58] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_99 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[57] WL[56] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_100 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[55] WL[54] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_101 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[53] WL[52] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_102 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[51] WL[50] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_103 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[49] WL[48] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_104 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[47] WL[46] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_105 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[45] WL[44] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_106 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[43] WL[42] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_107 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[41] WL[40] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_108 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[39] WL[38] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_109 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[37] WL[36] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_110 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[35] WL[34] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_111 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[33] WL[32] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_112 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[31] WL[30] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_113 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[29] WL[28] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_114 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[27] WL[26] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_115 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[25] WL[24] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_116 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[23] WL[22] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_117 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[21] WL[20] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_118 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[19] WL[18] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_119 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[17] WL[16] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_120 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[15] WL[14] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_121 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[13] WL[12] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_122 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[11] WL[10] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_123 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[9] WL[8] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_124 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[7] WL[6] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_125 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[5] WL[4] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_126 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[3] WL[2] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
XIS013EELPSP_127 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell2x2
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcellx4_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcellx4_b VDDC VSS WL[3] WL[2] WL[1] WL[0]
XIBITCELL_0 net016 net18 VDDC VSS WL[0] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_1 net27 net23 VDDC VSS WL[2] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_2 net016 net18 VDDC VSS WL[1] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_3 net27 net23 VDDC VSS WL[3] S013LLLPSP_X256Y8D8_BITCELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell4x2_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell4x2_b VDDC VSS WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 VDDC VSS WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcellx4_b
XIS013EELPSP_1 VDDC VSS WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcellx4_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] VDDC VSS S013LLLPSP_X256Y8D8_S013EELPSP_bitcellredundance2x2
XIS013EELPSP_1 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192]
+WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182]
+WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172]
+WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162]
+WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152]
+WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142]
+WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132]
+WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122]
+WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112]
+WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102]
+WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92]
+WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82]
+WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72]
+WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2
XIS013EELPSP_2 VDDC VSS STWL[3] STWL[2] STWL[1] STWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell4x2_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL B BX VDDC VSS WL
MM5 BCN BC VDDC VDDC PL W=160.000n L=150.00n m=1
MM6 BC BCN VDDC VDDC PL W=160.000n L=150.00n m=1
MM0 BCN BC VSS VSS NPD W=220.00n L=130.00n m=1
MM1 BC BCN VSS VSS NPD W=220.00n L=130.00n m=1
MM2 BX WL BCN VSS NPG W=150.000n L=175.00n m=1
MM3 B VSS BC VSS NPG W=150.000n L=175.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL_b STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS
XIS013EELPSP_0 net28 net19 VDDC VSS STWL[2] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL
XIS013EELPSP_1 net012 net14 VDDC VSS STWL[1] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL
XIBITCELL_2 net28 net19 VDDC VSS STWL[3] S013LLLPSP_X256Y8D8_BITCELL
XIBITCELL_3 net012 net14 VDDC VSS STWL[0] S013LLLPSP_X256Y8D8_BITCELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR_MID
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR_MID BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] VDDC VSS S013LLLPSP_X256Y8D8_S013EELPSP_bitcellredundance2x2
XIS013EELPSP_1 BL[1] BL[0] BLX[1] BLX[0] VDDC VSS WL[255] WL[254] WL[253] WL[252]
+WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242]
+WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232]
+WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222]
+WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212]
+WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202]
+WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192]
+WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182]
+WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172]
+WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162]
+WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152]
+WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142]
+WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132]
+WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122]
+WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112]
+WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102]
+WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92]
+WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82]
+WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72]
+WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62]
+WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52]
+WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42]
+WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32]
+WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22]
+WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2]
+WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2
XIS013EELPSP_2 VDDC VSS STWL[3] STWL[2] STWL[1] STWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcellx4_b
XIS013EELPSP_3 STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS S013LLLPSP_X256Y8D8_S013EELPSP_bitcell_STWL_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_MID_BW
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_MID_BW BWEN D DCTRCLK DCTRCLKX Q RWL[1] RWL[0] SACK1 SACK4 STWL[3]
+STWL[2] STWL[1] STWL[0] VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0]
XIS013EELPSP_0 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6]
+BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] BWEN DCTRCLK DCTRCLKX D
+Q SACK1 SACK4 VDDP VSS WE YX[7] YX[6] YX[5] YX[4]
+YX[3] YX[2] YX[1] YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMX8SAWR_BW
XIS013EELPSP_1 BL[7] BL[6] BLX[7] BLX[6] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_2 BL[5] BL[4] BLX[5] BLX[4] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_3 BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_4 BL[3] BL[2] BLX[3] BLX[2] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR_MID
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW BWEN D DCTRCLK DCTRCLKX Q RWL[1] RWL[0] SACK1 SACK4 STWL[3]
+STWL[2] STWL[1] STWL[0] VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0]
XIS013EELPSP_0 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6]
+BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] BWEN DCTRCLK DCTRCLKX D
+Q SACK1 SACK4 VDDP VSS WE YX[7] YX[6] YX[5] YX[4]
+YX[3] YX[2] YX[1] YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_YMX8SAWR_BW
XIS013EELPSP_1 BL[7] BL[6] BLX[7] BLX[6] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_2 BL[5] BL[4] BLX[5] BLX[4] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_3 BL[3] BL[2] BLX[3] BLX[2] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
XIS013EELPSP_4 BL[1] BL[0] BLX[1] BLX[0] RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0]
+VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_bitcell256x2abR
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_STRAP_CELL
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_STRAP_CELL WL VSS
MN0 VSS WL VSS VSS N15LL W=0.075u L=0.175u m=1
MN1 VSS WL VSS VSS N15LL W=0.075u L=0.175u m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_strap256
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_strap256 WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] VSS
XISTRAP_0 WL[0] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_1 WL[1] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_2 WL[2] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_3 WL[3] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_4 WL[4] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_5 WL[5] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_6 WL[6] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_7 WL[7] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_8 WL[8] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_9 WL[9] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_10 WL[10] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_11 WL[11] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_12 WL[12] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_13 WL[13] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_14 WL[14] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_15 WL[15] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_16 WL[16] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_17 WL[17] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_18 WL[18] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_19 WL[19] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_20 WL[20] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_21 WL[21] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_22 WL[22] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_23 WL[23] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_24 WL[24] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_25 WL[25] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_26 WL[26] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_27 WL[27] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_28 WL[28] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_29 WL[29] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_30 WL[30] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_31 WL[31] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_32 WL[32] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_33 WL[33] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_34 WL[34] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_35 WL[35] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_36 WL[36] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_37 WL[37] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_38 WL[38] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_39 WL[39] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_40 WL[40] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_41 WL[41] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_42 WL[42] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_43 WL[43] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_44 WL[44] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_45 WL[45] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_46 WL[46] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_47 WL[47] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_48 WL[48] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_49 WL[49] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_50 WL[50] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_51 WL[51] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_52 WL[52] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_53 WL[53] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_54 WL[54] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_55 WL[55] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_56 WL[56] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_57 WL[57] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_58 WL[58] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_59 WL[59] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_60 WL[60] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_61 WL[61] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_62 WL[62] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_63 WL[63] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_64 WL[64] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_65 WL[65] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_66 WL[66] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_67 WL[67] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_68 WL[68] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_69 WL[69] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_70 WL[70] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_71 WL[71] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_72 WL[72] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_73 WL[73] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_74 WL[74] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_75 WL[75] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_76 WL[76] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_77 WL[77] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_78 WL[78] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_79 WL[79] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_80 WL[80] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_81 WL[81] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_82 WL[82] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_83 WL[83] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_84 WL[84] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_85 WL[85] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_86 WL[86] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_87 WL[87] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_88 WL[88] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_89 WL[89] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_90 WL[90] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_91 WL[91] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_92 WL[92] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_93 WL[93] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_94 WL[94] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_95 WL[95] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_96 WL[96] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_97 WL[97] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_98 WL[98] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_99 WL[99] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_100 WL[100] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_101 WL[101] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_102 WL[102] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_103 WL[103] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_104 WL[104] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_105 WL[105] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_106 WL[106] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_107 WL[107] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_108 WL[108] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_109 WL[109] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_110 WL[110] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_111 WL[111] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_112 WL[112] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_113 WL[113] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_114 WL[114] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_115 WL[115] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_116 WL[116] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_117 WL[117] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_118 WL[118] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_119 WL[119] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_120 WL[120] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_121 WL[121] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_122 WL[122] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_123 WL[123] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_124 WL[124] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_125 WL[125] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_126 WL[126] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_127 WL[127] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_128 WL[128] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_129 WL[129] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_130 WL[130] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_131 WL[131] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_132 WL[132] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_133 WL[133] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_134 WL[134] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_135 WL[135] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_136 WL[136] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_137 WL[137] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_138 WL[138] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_139 WL[139] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_140 WL[140] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_141 WL[141] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_142 WL[142] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_143 WL[143] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_144 WL[144] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_145 WL[145] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_146 WL[146] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_147 WL[147] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_148 WL[148] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_149 WL[149] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_150 WL[150] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_151 WL[151] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_152 WL[152] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_153 WL[153] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_154 WL[154] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_155 WL[155] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_156 WL[156] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_157 WL[157] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_158 WL[158] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_159 WL[159] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_160 WL[160] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_161 WL[161] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_162 WL[162] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_163 WL[163] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_164 WL[164] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_165 WL[165] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_166 WL[166] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_167 WL[167] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_168 WL[168] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_169 WL[169] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_170 WL[170] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_171 WL[171] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_172 WL[172] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_173 WL[173] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_174 WL[174] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_175 WL[175] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_176 WL[176] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_177 WL[177] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_178 WL[178] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_179 WL[179] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_180 WL[180] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_181 WL[181] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_182 WL[182] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_183 WL[183] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_184 WL[184] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_185 WL[185] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_186 WL[186] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_187 WL[187] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_188 WL[188] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_189 WL[189] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_190 WL[190] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_191 WL[191] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_192 WL[192] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_193 WL[193] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_194 WL[194] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_195 WL[195] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_196 WL[196] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_197 WL[197] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_198 WL[198] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_199 WL[199] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_200 WL[200] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_201 WL[201] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_202 WL[202] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_203 WL[203] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_204 WL[204] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_205 WL[205] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_206 WL[206] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_207 WL[207] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_208 WL[208] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_209 WL[209] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_210 WL[210] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_211 WL[211] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_212 WL[212] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_213 WL[213] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_214 WL[214] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_215 WL[215] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_216 WL[216] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_217 WL[217] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_218 WL[218] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_219 WL[219] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_220 WL[220] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_221 WL[221] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_222 WL[222] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_223 WL[223] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_224 WL[224] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_225 WL[225] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_226 WL[226] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_227 WL[227] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_228 WL[228] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_229 WL[229] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_230 WL[230] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_231 WL[231] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_232 WL[232] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_233 WL[233] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_234 WL[234] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_235 WL[235] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_236 WL[236] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_237 WL[237] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_238 WL[238] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_239 WL[239] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_240 WL[240] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_241 WL[241] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_242 WL[242] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_243 WL[243] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_244 WL[244] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_245 WL[245] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_246 WL[246] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_247 WL[247] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_248 WL[248] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_249 WL[249] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_250 WL[250] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_251 WL[251] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_252 WL[252] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_253 WL[253] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_254 WL[254] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_255 WL[255] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_strap_STWL_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_strap_STWL_b STWL[3] STWL[2] STWL[1] STWL[0] VSS
XISTRAP_0 STWL[1] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_1 STWL[3] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_2 STWL[2] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_3 STWL[0] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0] VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0]
XISTRAP_0 RWL[1] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XISTRAP_1 RWL[0] VSS S013LLLPSP_X256Y8D8_STRAP_CELL
XIS013EELPSP_2 WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246]
+WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236]
+WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226]
+WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216]
+WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206]
+WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196]
+WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186]
+WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176]
+WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166]
+WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156]
+WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146]
+WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136]
+WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126]
+WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116]
+WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106]
+WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96]
+WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86]
+WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76]
+WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66]
+WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56]
+WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46]
+WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36]
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26]
+WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16]
+WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6]
+WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] VSS S013LLLPSP_X256Y8D8_S013EELPSP_strap256
XIS013EELPSP_3 STWL[3] STWL[2] STWL[1] STWL[0] VSS S013LLLPSP_X256Y8D8_S013EELPSP_strap_STWL_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap B BX VDDC VSS WL
MM2 BX WL net034 VSS NPG W=150.000n L=175.00n m=1
MTA1 B WL net27 VSS NPG W=150.000n L=175.00n m=1
MM1 net034 net27 VSS VSS NPD W=220.000n L=130.000n m=1
MTD1 net27 net034 VSS VSS NPD W=220.000n L=130.000n m=1
MM0 net034 net27 VDDC VDDC PL W=160.000n L=150.000n m=1
MTL1 net27 net034 VDDC VDDC PL W=160.000n L=150.000n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4 VDDC VSS WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 net28 net26 VDDC VSS WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_1 net28 net26 VDDC VSS WL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_2 net38 net36 VDDC VSS WL[2] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_3 net38 net36 VDDC VSS WL[3] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap256
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap256 VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 VDDC VSS WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_1 VDDC VSS WL[7] WL[6] WL[5] WL[4] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_2 VDDC VSS WL[11] WL[10] WL[9] WL[8] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_3 VDDC VSS WL[15] WL[14] WL[13] WL[12] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_4 VDDC VSS WL[19] WL[18] WL[17] WL[16] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_5 VDDC VSS WL[23] WL[22] WL[21] WL[20] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_6 VDDC VSS WL[27] WL[26] WL[25] WL[24] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_7 VDDC VSS WL[31] WL[30] WL[29] WL[28] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_8 VDDC VSS WL[35] WL[34] WL[33] WL[32] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_9 VDDC VSS WL[39] WL[38] WL[37] WL[36] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_10 VDDC VSS WL[43] WL[42] WL[41] WL[40] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_11 VDDC VSS WL[47] WL[46] WL[45] WL[44] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_12 VDDC VSS WL[51] WL[50] WL[49] WL[48] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_13 VDDC VSS WL[55] WL[54] WL[53] WL[52] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_14 VDDC VSS WL[59] WL[58] WL[57] WL[56] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_15 VDDC VSS WL[63] WL[62] WL[61] WL[60] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_16 VDDC VSS WL[67] WL[66] WL[65] WL[64] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_17 VDDC VSS WL[71] WL[70] WL[69] WL[68] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_18 VDDC VSS WL[75] WL[74] WL[73] WL[72] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_19 VDDC VSS WL[79] WL[78] WL[77] WL[76] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_20 VDDC VSS WL[83] WL[82] WL[81] WL[80] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_21 VDDC VSS WL[87] WL[86] WL[85] WL[84] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_22 VDDC VSS WL[91] WL[90] WL[89] WL[88] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_23 VDDC VSS WL[95] WL[94] WL[93] WL[92] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_24 VDDC VSS WL[99] WL[98] WL[97] WL[96] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_25 VDDC VSS WL[103] WL[102] WL[101] WL[100] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_26 VDDC VSS WL[107] WL[106] WL[105] WL[104] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_27 VDDC VSS WL[111] WL[110] WL[109] WL[108] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_28 VDDC VSS WL[115] WL[114] WL[113] WL[112] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_29 VDDC VSS WL[119] WL[118] WL[117] WL[116] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_30 VDDC VSS WL[123] WL[122] WL[121] WL[120] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_31 VDDC VSS WL[127] WL[126] WL[125] WL[124] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_32 VDDC VSS WL[131] WL[130] WL[129] WL[128] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_33 VDDC VSS WL[135] WL[134] WL[133] WL[132] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_34 VDDC VSS WL[139] WL[138] WL[137] WL[136] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_35 VDDC VSS WL[143] WL[142] WL[141] WL[140] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_36 VDDC VSS WL[147] WL[146] WL[145] WL[144] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_37 VDDC VSS WL[151] WL[150] WL[149] WL[148] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_38 VDDC VSS WL[155] WL[154] WL[153] WL[152] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_39 VDDC VSS WL[159] WL[158] WL[157] WL[156] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_40 VDDC VSS WL[163] WL[162] WL[161] WL[160] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_41 VDDC VSS WL[167] WL[166] WL[165] WL[164] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_42 VDDC VSS WL[171] WL[170] WL[169] WL[168] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_43 VDDC VSS WL[175] WL[174] WL[173] WL[172] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_44 VDDC VSS WL[179] WL[178] WL[177] WL[176] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_45 VDDC VSS WL[183] WL[182] WL[181] WL[180] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_46 VDDC VSS WL[187] WL[186] WL[185] WL[184] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_47 VDDC VSS WL[191] WL[190] WL[189] WL[188] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_48 VDDC VSS WL[195] WL[194] WL[193] WL[192] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_49 VDDC VSS WL[199] WL[198] WL[197] WL[196] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_50 VDDC VSS WL[203] WL[202] WL[201] WL[200] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_51 VDDC VSS WL[207] WL[206] WL[205] WL[204] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_52 VDDC VSS WL[211] WL[210] WL[209] WL[208] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_53 VDDC VSS WL[215] WL[214] WL[213] WL[212] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_54 VDDC VSS WL[219] WL[218] WL[217] WL[216] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_55 VDDC VSS WL[223] WL[222] WL[221] WL[220] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_56 VDDC VSS WL[227] WL[226] WL[225] WL[224] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_57 VDDC VSS WL[231] WL[230] WL[229] WL[228] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_58 VDDC VSS WL[235] WL[234] WL[233] WL[232] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_59 VDDC VSS WL[239] WL[238] WL[237] WL[236] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_60 VDDC VSS WL[243] WL[242] WL[241] WL[240] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_61 VDDC VSS WL[247] WL[246] WL[245] WL[244] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_62 VDDC VSS WL[251] WL[250] WL[249] WL[248] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
XIS013EELPSP_63 VDDC VSS WL[255] WL[254] WL[253] WL[252] S013LLLPSP_X256Y8D8_S013EELPSP_pcapx4
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_b STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS
XIS013EELPSP_0 net029 net027 VDDC VSS STWL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_1 net14 net019 VDDC VSS STWL[3] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_2 net14 net019 VDDC VSS STWL[2] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_3 net029 net027 VDDC VSS STWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge256
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge256 RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 net031 net25 VDDC VSS RWL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_1 net031 net25 VDDC VSS RWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap
XIS013EELPSP_2 VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap256
XIS013EELPSP_3 STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st B BX VDDC VSS WL0
MTL1 net42 net51 VDDC VDDC PL W=160.000n L=150.000n m=1
MTL0 net51 net42 VDDC VDDC PL W=160.000n L=150.000n m=1
MTD0 net51 net42 VSS VSS NPD W=220.000n L=130.000n m=1
MTD1 net42 net51 VSS VSS NPD W=220.000n L=130.000n m=1
MTA0 B WL0 net51 VSS NPG W=150.000n L=175.00n m=1
MTA1 BX VSS net42 VSS NPG W=150.000n L=175.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4 BX VDDC VSS WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 net32 BX VDDC VSS WL[3] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_1 net32 BX VDDC VSS WL[2] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_2 net42 BX VDDC VSS WL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_3 net42 BX VDDC VSS WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st256
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st256 BX VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249]
+WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239]
+WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229]
+WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219]
+WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209]
+WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199]
+WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189]
+WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179]
+WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169]
+WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159]
+WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149]
+WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139]
+WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129]
+WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119]
+WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109]
+WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99]
+WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89]
+WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79]
+WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69]
+WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 BX VDDC VSS WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_1 BX VDDC VSS WL[7] WL[6] WL[5] WL[4] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_2 BX VDDC VSS WL[11] WL[10] WL[9] WL[8] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_3 BX VDDC VSS WL[15] WL[14] WL[13] WL[12] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_4 BX VDDC VSS WL[19] WL[18] WL[17] WL[16] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_5 BX VDDC VSS WL[23] WL[22] WL[21] WL[20] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_6 BX VDDC VSS WL[27] WL[26] WL[25] WL[24] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_7 BX VDDC VSS WL[31] WL[30] WL[29] WL[28] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_8 BX VDDC VSS WL[35] WL[34] WL[33] WL[32] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_9 BX VDDC VSS WL[39] WL[38] WL[37] WL[36] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_10 BX VDDC VSS WL[43] WL[42] WL[41] WL[40] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_11 BX VDDC VSS WL[47] WL[46] WL[45] WL[44] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_12 BX VDDC VSS WL[51] WL[50] WL[49] WL[48] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_13 BX VDDC VSS WL[55] WL[54] WL[53] WL[52] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_14 BX VDDC VSS WL[59] WL[58] WL[57] WL[56] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_15 BX VDDC VSS WL[63] WL[62] WL[61] WL[60] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_16 BX VDDC VSS WL[67] WL[66] WL[65] WL[64] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_17 BX VDDC VSS WL[71] WL[70] WL[69] WL[68] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_18 BX VDDC VSS WL[75] WL[74] WL[73] WL[72] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_19 BX VDDC VSS WL[79] WL[78] WL[77] WL[76] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_20 BX VDDC VSS WL[83] WL[82] WL[81] WL[80] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_21 BX VDDC VSS WL[87] WL[86] WL[85] WL[84] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_22 BX VDDC VSS WL[91] WL[90] WL[89] WL[88] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_23 BX VDDC VSS WL[95] WL[94] WL[93] WL[92] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_24 BX VDDC VSS WL[99] WL[98] WL[97] WL[96] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_25 BX VDDC VSS WL[103] WL[102] WL[101] WL[100] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_26 BX VDDC VSS WL[107] WL[106] WL[105] WL[104] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_27 BX VDDC VSS WL[111] WL[110] WL[109] WL[108] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_28 BX VDDC VSS WL[115] WL[114] WL[113] WL[112] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_29 BX VDDC VSS WL[119] WL[118] WL[117] WL[116] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_30 BX VDDC VSS WL[123] WL[122] WL[121] WL[120] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_31 BX VDDC VSS WL[127] WL[126] WL[125] WL[124] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_32 BX VDDC VSS WL[131] WL[130] WL[129] WL[128] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_33 BX VDDC VSS WL[135] WL[134] WL[133] WL[132] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_34 BX VDDC VSS WL[139] WL[138] WL[137] WL[136] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_35 BX VDDC VSS WL[143] WL[142] WL[141] WL[140] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_36 BX VDDC VSS WL[147] WL[146] WL[145] WL[144] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_37 BX VDDC VSS WL[151] WL[150] WL[149] WL[148] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_38 BX VDDC VSS WL[155] WL[154] WL[153] WL[152] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_39 BX VDDC VSS WL[159] WL[158] WL[157] WL[156] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_40 BX VDDC VSS WL[163] WL[162] WL[161] WL[160] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_41 BX VDDC VSS WL[167] WL[166] WL[165] WL[164] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_42 BX VDDC VSS WL[171] WL[170] WL[169] WL[168] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_43 BX VDDC VSS WL[175] WL[174] WL[173] WL[172] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_44 BX VDDC VSS WL[179] WL[178] WL[177] WL[176] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_45 BX VDDC VSS WL[183] WL[182] WL[181] WL[180] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_46 BX VDDC VSS WL[187] WL[186] WL[185] WL[184] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_47 BX VDDC VSS WL[191] WL[190] WL[189] WL[188] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_48 BX VDDC VSS WL[195] WL[194] WL[193] WL[192] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_49 BX VDDC VSS WL[199] WL[198] WL[197] WL[196] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_50 BX VDDC VSS WL[203] WL[202] WL[201] WL[200] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_51 BX VDDC VSS WL[207] WL[206] WL[205] WL[204] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_52 BX VDDC VSS WL[211] WL[210] WL[209] WL[208] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_53 BX VDDC VSS WL[215] WL[214] WL[213] WL[212] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_54 BX VDDC VSS WL[219] WL[218] WL[217] WL[216] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_55 BX VDDC VSS WL[223] WL[222] WL[221] WL[220] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_56 BX VDDC VSS WL[227] WL[226] WL[225] WL[224] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_57 BX VDDC VSS WL[231] WL[230] WL[229] WL[228] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_58 BX VDDC VSS WL[235] WL[234] WL[233] WL[232] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_59 BX VDDC VSS WL[239] WL[238] WL[237] WL[236] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_60 BX VDDC VSS WL[243] WL[242] WL[241] WL[240] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_61 BX VDDC VSS WL[247] WL[246] WL[245] WL[244] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_62 BX VDDC VSS WL[251] WL[250] WL[249] WL[248] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
XIS013EELPSP_63 BX VDDC VSS WL[255] WL[254] WL[253] WL[252] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_stx4
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_st_b
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_st_b STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS
XIS013EELPSP_0 net14 net28 VDDC VSS STWL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_1 net24 net18 VDDC VSS STWL[3] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_2 net24 net18 VDDC VSS STWL[2] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_3 net14 net28 VDDC VSS STWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge_st256
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge_st256 BL RWL[1] RWL[0] STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0]
XIS013EELPSP_0 net031 BL VDDC VSS RWL[1] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_1 net031 BL VDDC VSS RWL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st
XIS013EELPSP_2 BL VDDC VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249]
+WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239]
+WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229]
+WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219]
+WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209]
+WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199]
+WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189]
+WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179]
+WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169]
+WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159]
+WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149]
+WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139]
+WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129]
+WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119]
+WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109]
+WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99]
+WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89]
+WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79]
+WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69]
+WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59]
+WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39]
+WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29]
+WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19]
+WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_st256
XIS013EELPSP_3 STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS S013LLLPSP_X256Y8D8_S013EELPSP_pcap_STWL_st_b
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_right
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_right BWEN[3] BWEN[2] BWEN[1] BWEN[0] D[3] D[2] D[1] D[0] DBL DCTRCLK
+DCTRCLKX Q[3] Q[2] Q[1] Q[0] RWL[1] RWL[0] SACK1 SACK4 STWL
+VDDP VDDC VSS WE WL[255] WL[254] WL[253] WL[252] WL[251] WL[250]
+WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240]
+WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230]
+WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220]
+WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210]
+WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200]
+WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190]
+WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180]
+WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170]
+WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160]
+WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150]
+WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140]
+WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130]
+WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120]
+WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110]
+WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100]
+WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90]
+WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80]
+WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70]
+WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60]
+WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50]
+WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40]
+WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30]
+WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20]
+WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10]
+WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
+YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0]
XIS013EELPSP_0 BWEN[2] D[2] DCTRCLK DCTRCLKX Q[2] RWL[1] RWL[0] SACK1 SACK4 VSS
+STWL STWL VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_MID_BW
XIS013EELPSP_1 BWEN[0] D[0] DCTRCLK DCTRCLKX Q[0] RWL[1] RWL[0] SACK1 SACK4 VSS
+STWL STWL VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_2 BWEN[1] D[1] DCTRCLK DCTRCLKX Q[1] RWL[1] RWL[0] SACK1 SACK4 VSS
+STWL STWL VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_3 BWEN[3] D[3] DCTRCLK DCTRCLKX Q[3] RWL[1] RWL[0] SACK1 SACK4 VSS
+VSS VSS VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_4 RWL[1] RWL[0] VSS STWL STWL VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_5 RWL[1] RWL[0] VSS STWL STWL VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_6 RWL[1] RWL[0] VSS VSS VSS VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_7 RWL[1] RWL[0] VSS VSS VSS VSS VDDC VSS WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge256
XIS013EELPSP_8 DBL RWL[1] RWL[0] VSS STWL STWL VSS VDDC VSS WL[255]
+WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245]
+WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235]
+WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215]
+WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205]
+WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195]
+WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175]
+WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165]
+WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155]
+WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135]
+WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125]
+WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115]
+WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95]
+WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85]
+WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75]
+WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55]
+WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45]
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35]
+WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15]
+WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5]
+WL[4] WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge_st256
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_left
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_left BWEN[3] BWEN[2] BWEN[1] BWEN[0] D[3] D[2] D[1] D[0] DCTRCLK DCTRCLKX
+Q[3] Q[2] Q[1] Q[0] RWLU[1] RWLU[0] SACK1 SACK4 VDDP VDDC
+VSS WE WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248]
+WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238]
+WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228]
+WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218]
+WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208]
+WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] WL[198]
+WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] WL[189] WL[188]
+WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178]
+WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168]
+WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158]
+WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148]
+WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138]
+WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128]
+WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118]
+WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] WL[108]
+WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] WL[99] WL[98]
+WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] WL[88]
+WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78]
+WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68]
+WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58]
+WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48]
+WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38]
+WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28]
+WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18]
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8]
+WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0]
XIS013EELPSP_0 BWEN[0] D[0] DCTRCLK DCTRCLKX Q[0] RWLU[1] RWLU[0] SACK1 SACK4 VSS
+VSS VSS VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_1 BWEN[1] D[1] DCTRCLK DCTRCLKX Q[1] RWLU[1] RWLU[0] SACK1 SACK4 VSS
+VSS VSS VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_2 BWEN[2] D[2] DCTRCLK DCTRCLKX Q[2] RWLU[1] RWLU[0] SACK1 SACK4 VSS
+VSS VSS VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_3 BWEN[3] D[3] DCTRCLK DCTRCLKX Q[3] RWLU[1] RWLU[0] SACK1 SACK4 VSS
+VSS VSS VSS VDDP VDDC VSS WE WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1]
+YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D1_BW
XIS013EELPSP_4 RWLU[1] RWLU[0] VSS VSS VSS VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_5 RWLU[1] RWLU[0] VSS VSS VSS VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_6 RWLU[1] RWLU[0] VSS VSS VSS VSS VSS WL[255] WL[254] WL[253]
+WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] WL[243]
+WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223]
+WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213]
+WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203]
+WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183]
+WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173]
+WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163]
+WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144] WL[143]
+WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133]
+WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123]
+WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103]
+WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93]
+WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83]
+WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63]
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53]
+WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43]
+WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23]
+WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13]
+WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3]
+WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_X256_Y8_strap
XIS013EELPSP_7 RWLU[1] RWLU[0] VSS VSS VSS VSS VDDC VSS WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge256
XIS013EELPSP_8 RWLU[1] RWLU[0] VSS VSS VSS VSS VDDC VSS WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0] S013LLLPSP_X256Y8D8_S013EELPSP_pcap_edge256
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_left
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_left CLK CLKX RDE RWLL VDDP VSS WLCKX
MP9 net64 net97 VDDP VDDP P15LL W=4u L=130.00n m=1
XI114 net64 net97 net93 VDDP VSS WLCKX / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI2 net73 CLKX CLK VDDP VSS net69 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI3 net77 VDDP VSS net73 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI8 RDE VDDP VSS net77 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI129 net64 VDDP VSS RWLL / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=2u
XI1 net93 VDDP VSS net69 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI0 net69 VDDP VSS net93 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI24 net93 VDDP VSS net97 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_right
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_right CLK CLKX RDE RWLR VDDP VSS WLCKX
MP0 net58 net97 VDDP VDDP P15LL W=4u L=130.00n m=1
XI5 net58 net97 net93 VDDP VSS WLCKX / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI2 net73 CLKX CLK VDDP VSS net69 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI3 net77 VDDP VSS net73 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI8 RDE VDDP VSS net77 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI7 net58 VDDP VSS RWLR / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=2u
XI1 net93 VDDP VSS net69 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI0 net69 VDDP VSS net93 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI24 net93 VDDP VSS net97 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_STWL_DEC
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_STWL_DEC EMCLK STWL VDDP VSS
MP9 A T_HIGH VDDP VDDP P15LL W=800.0n L=130.00n m=1
MP18 net61 net61 VDDP VDDP P15LL W=800.0n L=130.00n m=1
MM4 T_HIGH net77 VDDP VDDP P15LL W=2u L=130.00n m=1
MM0 STWL C VDDP VDDP P15LL W=5u L=130.00n m=1
MM5 net77 net77 VSS VSS N15LL W=800.0n L=130.00n m=1
MN18 T_LOW net61 VSS VSS N15LL W=1u L=130.00n m=1
MM1 STWL C VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS C / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=3u nl=130.00n nw=3u
XI8 A VDDP VSS B / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1u nl=130.00n nw=1u
XI114 A T_HIGH T_LOW VDDP VSS EMCLK / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=800.0n nl=130.00n  nw=1.2u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH_S
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH_S Tie_high VDDP VSS
MN18 net15 net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 Tie_high net15 VDDP VDDP P15LL W=3u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_nor2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_nor2 A B VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
MM3 Y B VSS VSS N15LL W=nw L=nl m=1
MM2 Y A VSS VSS N15LL W=nw L=nl m=1
MM1 Y B net35 VDDP P15LL W=pw L=pl m=1
MM0 net35 A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_OPDEC
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_OPDEC OP[1] OP[0] S[2] S[1] S[0] VDDP VSS
XI12 AX BX VDDP VSS S[2] / S013LLLPSP_X256Y8D8_nor2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI6 AX BX VDDP VSS S[0] / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI7 BX VDDP VSS S[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI1 OP[1] VDDP VSS BX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI0 OP[0] VDDP VSS AX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DischargeCells
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DischargeCells DUM_BL EMCLK S[2] S[1] S[0] VDDP VSS
MN6 net30 S[2] VSS VSS NPD W=220.000n L=130.000n m=8
MN5 net34 S[1] VSS VSS NPD W=220.000n L=130.000n m=4
MN2 net38 S[0] VSS VSS NPD W=220.000n L=130.000n m=4
MN1 net42 VDDP VSS VSS NPD W=220.000n L=130.000n m=4
MN16 DUM_BL EMCLK net42 VSS NPG W=150.000n L=175.00n m=4
MN7 DUM_BL EMCLK net30 VSS NPG W=150.000n L=175.00n m=8
MN4 DUM_BL EMCLK net34 VSS NPG W=150.000n L=175.00n m=4
MN3 DUM_BL EMCLK net38 VSS NPG W=150.000n L=175.00n m=4
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL_S
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL_S TieL VDDP VSS
MN18 TieL net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 net15 net15 VDDP VDDP P15LL W=1.6u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_SOP01
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_SOP01 DBL_right EMCLK STWL_right VDDP VSS
XI16 TieLS VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH_S
MM0 TieHS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 TieLS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 TieHS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 TieLS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_DischargeCells
XI21 TieLS TieHS OP[2] OP[1] OP[0] VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_OPDEC
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_ESDA14
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_ESDA14 A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2]
+A[1] A[0] CEN CLK S[1] S[0] VDDP VSS WEN
MM0 A[10] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM1110 A[11] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN29 A[5] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN30 A[6] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN31 A[8] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN32 A[7] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM1 A[9] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN28 WEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 S[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM13 S[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN7 A[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN6 A[2] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN5 A[4] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN4 A[3] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 CEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN2 A[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN0 CLK VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP29 A[5] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP30 A[6] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP31 A[8] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP32 A[7] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP28 WEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM2 A[10] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1112 A[11] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM3 A[9] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 S[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM15 S[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP7 A[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP6 A[2] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP5 A[4] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP4 A[3] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 CEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP2 A[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP0 CLK VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4 A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDDP VSS
XI19 net94 CLKX CLK VDDP VSS net70 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI18 net99 CLKX CLK VDDP VSS net76 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI14 net104 CLKX CLK VDDP VSS net82 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI10 net109 CLKX CLK VDDP VSS net88 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI21 AinX[0] Ain[1] VDDP VSS net94 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI20 Ain[0] Ain[1] VDDP VSS net99 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI15 Ain[0] AinX[1] VDDP VSS net104 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI9 AinX[0] AinX[1] VDDP VSS net109 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI25 net70 VDDP VSS PX[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI24 PX[2] VDDP VSS net70 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 PX[3] VDDP VSS net76 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI22 net76 VDDP VSS PX[3] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI17 net82 VDDP VSS PX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI16 PX[1] VDDP VSS net82 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI12 PX[0] VDDP VSS net88 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI11 net88 VDDP VSS PX[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI3 AinX[1] VDDP VSS Ain[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI2 A[1] VDDP VSS AinX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI1 AinX[0] VDDP VSS Ain[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI0 A[0] VDDP VSS AinX[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1.4u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PXA
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PXA A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] RDE VDDP VSS
XI19 net83 CLKX CLK VDDP VSS net59 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI18 net88 CLKX CLK VDDP VSS net65 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI14 net93 CLKX CLK VDDP VSS net71 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI10 net98 CLKX CLK VDDP VSS ALATCH / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI21 AinX[0] Ain[1] VDDP VSS net83 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI20 Ain[0] Ain[1] VDDP VSS net88 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI15 Ain[0] AinX[1] VDDP VSS net93 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI9 AinX[0] AinX[1] VDDP VSS net98 / S013LLLPSP_X256Y8D8_nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI62 A[0] VDDP VSS net100 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI25 net59 VDDP VSS PX[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI24 PX[2] VDDP VSS net59 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 PX[3] VDDP VSS net65 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI22 net65 VDDP VSS PX[3] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI17 net71 VDDP VSS PX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI16 PX[1] VDDP VSS net71 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI12 PX[0] VDDP VSS ALATCH / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI11 ALATCH VDDP VSS PX[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=7u nl=130.00n nw=2u
XI3 AinX[1] VDDP VSS Ain[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI2 A[1] VDDP VSS AinX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI1 net100 RDE VDDP VSS Ain[0] / S013LLLPSP_X256Y8D8_nor2 pl=130.00n pw=2u nl=130.00n nw=1u
XI0 A[0] RDE VDDP VSS AinX[0] / S013LLLPSP_X256Y8D8_nor2 pl=130.00n pw=1.5u nl=130.00n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_nand3
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_nand3 A B C VDDP VSS Y pw=1u pl=180.0n nw=1u nl=180.0n
MM6 net29 C VSS VSS N15LL W=nw L=nl m=1
MM5 net33 B net29 VSS N15LL W=nw L=nl m=1
MM4 Y A net33 VSS N15LL W=nw L=nl m=1
MM3 Y A VDDP VDDP P15LL W=pw L=pl m=1
MM2 Y B VDDP VDDP P15LL W=pw L=pl m=1
MM1 Y C VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC A[0] A[1] A[2] CLK CLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] VDDP VSS WLCKX
XI191 net270 WLCKX VDDP VSS net135 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI192 net326 WLCKX VDDP VSS net140 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI185 net274 WLCKX VDDP VSS net145 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI203 net286 WLCKX VDDP VSS net150 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI204 net282 WLCKX VDDP VSS net155 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI205 net318 WLCKX VDDP VSS net160 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI206 net278 WLCKX VDDP VSS net165 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI183 net314 WLCKX VDDP VSS net170 / S013LLLPSP_X256Y8D8_nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI186 net221 CLKX CLK VDDP VSS net175 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI194 net227 CLKX CLK VDDP VSS net181 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI193 net233 CLKX CLK VDDP VSS net187 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI207 net239 CLKX CLK VDDP VSS net193 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI208 net245 CLKX CLK VDDP VSS net199 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI209 net257 CLKX CLK VDDP VSS net205 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI210 net251 CLKX CLK VDDP VSS net211 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI134 net268 CLKX CLK VDDP VSS net0730 / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI187 Ain[0] AinX[1] AinX[2] VDDP VSS net221 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI196 AinX[0] Ain[1] AinX[2] VDDP VSS net227 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI195 Ain[0] Ain[1] AinX[2] VDDP VSS net233 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI211 AinX[0] Ain[1] Ain[2] VDDP VSS net239 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI212 Ain[0] Ain[1] Ain[2] VDDP VSS net245 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI214 AinX[0] AinX[1] Ain[2] VDDP VSS net251 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI213 Ain[0] AinX[1] Ain[2] VDDP VSS net257 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI133 AinX[0] AinX[1] AinX[2] VDDP VSS net268 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI229 net0346 VDDP VSS net270 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI228 net0334 VDDP VSS net274 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI234 net0182 VDDP VSS net278 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI232 net0370 VDDP VSS net282 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI231 net0277 VDDP VSS net286 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI188 net145 VDDP VSS FCKX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI189 net0334 VDDP VSS net175 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI237 A[2] VDDP VSS net298 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI235 A[0] VDDP VSS net302 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI199 net135 VDDP VSS FCKX[3] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI201 net0318 VDDP VSS net181 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI227 net359 VDDP VSS net314 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI233 net0342 VDDP VSS net318 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI220 net199 VDDP VSS net0370 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI230 net0318 VDDP VSS net326 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI82 net298 VDDP VSS Ain[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI215 net193 VDDP VSS net0277 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI217 net150 VDDP VSS FCKX[6] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI216 net0277 VDDP VSS net193 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI218 net155 VDDP VSS FCKX[7] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI138 Ain[2] VDDP VSS AinX[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI136 net359 VDDP VSS net0730 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI135 net0730 VDDP VSS net359 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI219 net0370 VDDP VSS net199 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI197 net187 VDDP VSS net0346 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI221 net205 VDDP VSS net0342 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI223 net160 VDDP VSS FCKX[5] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI224 net165 VDDP VSS FCKX[4] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI184 net170 VDDP VSS FCKX[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI225 net0182 VDDP VSS net211 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI190 net175 VDDP VSS net0334 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI222 net0342 VDDP VSS net205 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI226 net211 VDDP VSS net0182 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI198 net0346 VDDP VSS net187 / S013LLLPSP_X256Y8D8_inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI200 net140 VDDP VSS FCKX[2] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=5u nl=130.00n nw=5u
XI202 net181 VDDP VSS net0318 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI236 A[1] VDDP VSS net414 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI137 Ain[1] VDDP VSS AinX[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI2 net414 VDDP VSS Ain[1] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI132 Ain[0] VDDP VSS AinX[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
XI0 net302 VDDP VSS Ain[0] / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_OPDEC
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_OPDEC OP[1] OP[0] S[3] S[2] S[1] S[0] VDDP VSS
XI34 A BX VDDP VSS S[2] / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI35 A B VDDP VSS S[0] / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI27 AX BX VDDP VSS S[3] / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI31 AX B VDDP VSS S[1] / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI33 BX VDDP VSS B / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI32 AX VDDP VSS A / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI1 OP[1] VDDP VSS BX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI0 OP[0] VDDP VSS AX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_delay100p
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_delay100p VDDP VSS in out
MM0 net17 in VSS VSS N15LL W=800.0n L=300.00n m=1
MM1 net17 in VDDP VDDP P15LL W=800.0n L=130.00n m=1
XI0 net17 VDDP VSS out / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FIXDL
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FIXDL EMCLK IN OP[1] OP[0] VDDP VSS prc
XI22 VDDP VSS net36 net37 / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_delay100p
XI20 VDDP VSS net40 net36 / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_delay100p
XI19 VDDP VSS net44 net40 / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_delay100p
XI25 net37 SX[3] S[3] VDDP VSS EMCLK / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI126 net40 SX[1] S[1] VDDP VSS EMCLK / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI24 net36 SX[2] S[2] VDDP VSS EMCLK / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI144 net44 SX[0] S[0] VDDP VSS EMCLK / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=4u nl=130.00n nw=4u
XI136 IN VDDP VSS prc / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
XI137 prc VDDP VSS net44 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
XI3[3] S[3] VDDP VSS SX[3] / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[2] S[2] VDDP VSS SX[2] / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[1] S[1] VDDP VSS SX[1] / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[0] S[0] VDDP VSS SX[0] / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI0 OP[1] OP[0] S[3] S[2] S[1] S[0] VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_OPDEC
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_MUX2
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_MUX2 I0 I1 S VDDP VSS Z
XI2 net40 net44 VDDP VSS net030 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=2u nl=130n nw=1u
XI8 net030 VDDP VSS Z / S013LLLPSP_X256Y8D8_inv pl=130n pw=4u nl=130n nw=2u
XI6 net49 VDDP VSS net40 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2u nl=130n nw=1u
XI4 net54 VDDP VSS net44 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2u nl=130n nw=1u
XI5 S VDDP VSS net36 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2u nl=130n nw=1u
XI3 I0 net36 VDDP VSS net54 / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=2u nl=130.0n nw=1u
XI7 I1 S VDDP VSS net49 / S013LLLPSP_X256Y8D8_nand2 pl=130.0n pw=2u nl=130.0n nw=1u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_delayline_2p4
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_delayline_2p4 VDDP VSS Vin Vout
XI275 Vin VDDP VSS net145 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=1u
MM0 Vout net145 VDDP VDDP P15LL W=4u L=130.00n m=1
MM1 Vout net145 VSS VSS N15LL W=2u L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_buffer_split_right0_mode
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_buffer_split_right0_mode A SM VDDP VSS Y
XI143 A net0861 SM VDDP VSS Y / S013LLLPSP_X256Y8D8_MUX2
XI142 VDDP VSS A net0861 / S013LLLPSP_X256Y8D8_S013EELPSP_delayline_2p4
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_CLKDRV_mode_V1
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_CLKDRV_mode_V1 ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right DCTRCLK_right
+EMCLK FB_right INTCLKX INTCLKX_right S[1] S[0] SACK1 SACK1_right SACK4 SACK4_right
+SM VDDP VMINE VSS WE WEN WE_right
XI215 WE SM VDDP VSS WE_right / S013LLLPSP_X256Y8D8_buffer_split_right0_mode
XI197 CLKLATCH SM VDDP VSS net0257 / S013LLLPSP_X256Y8D8_buffer_split_right0_mode
XI173 EMCLK CLKLATCH S[1] S[0] VDDP VSS prc_right / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FIXDL
XI134 TESTB net285 VDDP VSS net168 / S013LLLPSP_X256Y8D8_nand2 pl=130n pw=3u nl=130n nw=3u
XI175 net0397 net0411 VDDP VSS net0194 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=6u nl=130n nw=3u
XI174 net0342 net0397 VDDP VSS net0199 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=5u nl=130n nw=5u
XI128 CENINT CLK_BUF VDDP VSS net173 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=2u nl=130n nw=1.0u
XI143 net337 PRESACK1 VDDP VSS net178 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=5u nl=130n nw=5u
XI151 PRESACK1 CLKD VDDP VSS net183 / S013LLLPSP_X256Y8D8_nor2 pl=130n pw=6u nl=130n nw=3u
MM2 net186 CEN net190 VSS N15LL W=2u L=130.00n m=1
MM3 net190 net261 VSS VSS N15LL W=2u L=130.00n m=1
MM5 CLKLATCH CLK_BUF net198 VSS N15LL W=20u L=130.00n m=1
MM6 net198 net0214 VSS VSS N15LL W=20u L=130.00n m=1
MM1 net186 CEN net205 VDDP P15LL W=2u L=130.00n m=1
MM0 net205 CLK_BUF VDDP VDDP P15LL W=2u L=130.00n m=1
MM11 CLKLATCH CLK_BUF up2 VDDP P15LL W=8.0u L=130.00n m=1
MM4 CLKLATCH net168 VDDP VDDP P15LL W=10u L=130.00n m=1
MM7 FB_right prc_right VDDP VDDP P15LL W=4.8u L=130.00n m=1
MM10 up2 TESTB VDDP VDDP P15LL W=8.0u L=130.00n m=1
XI114 net241 ACTRCLKX ACTRCLK VDDP VSS WENLATCH / S013LLLPSP_X256Y8D8_tgate pl=130n pw=2u nl=130n  nw=2u
XI212 net0397 VDDP VSS net0344 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI214 net0352 VDDP VSS net0227 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI209 CLK VDDP VSS net0222 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2.0000u nl=130n nw=1.2u
XI210 net0222 VDDP VSS CLK_BUF / S013LLLPSP_X256Y8D8_inv pl=130n pw=4u nl=130n nw=2.4u
XI169 VMINE VDDP VSS TESTB / S013LLLPSP_X256Y8D8_inv pl=130n pw=2.0u nl=130n nw=1.0u
XI188 net0397 VDDP VSS INTCLKX_right / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=10u
XI186 net0194 VDDP VSS SACK4_right / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=5u
XI177 net0257 VDDP VSS net0397 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=20u nl=130.00n nw=10u
XI183 net0199 VDDP VSS DCTRCLK_right / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI182 net0199 VDDP VSS net0326 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=6u nl=130.00n nw=6u
XI184 net0348 VDDP VSS net0330 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI179 net0199 VDDP VSS ACTRCLK_right / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI178 net0397 VDDP VSS net0257 / S013LLLPSP_X256Y8D8_inv pl=200.0n pw=250.00n nl=1u nw=250.00n
XI189 net0350 VDDP VSS net0342 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI185 net0330 VDDP VSS net0411 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI176 net0397 VDDP VSS net0350 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI181 net0326 VDDP VSS DCTRCLKX_right / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI180 ACTRCLK_right VDDP VSS ACTRCLKX_right / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n  nw=5u
XI110 WEN VDDP VSS net237 / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI211 net0344 VDDP VSS net0348 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI112 net237 VDDP VSS net241 / S013LLLPSP_X256Y8D8_inv pl=300n pw=2u nl=300n nw=2u
XI115 WENLATCH VDDP VSS net245 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2u nl=130n nw=2u
XI116 net245 VDDP VSS WENLATCH / S013LLLPSP_X256Y8D8_inv pl=300n pw=250.00n nl=600n nw=250.00n
XI208 net281 VDDP VSS net0214 / S013LLLPSP_X256Y8D8_inv pl=130n pw=6u nl=130n nw=3u
XI117 net245 VDDP VSS net253 / S013LLLPSP_X256Y8D8_inv pl=130n pw=6u nl=130n nw=4u
XI118 net253 VDDP VSS WE / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=5u
XI125 CLK_BUF VDDP VSS net261 / S013LLLPSP_X256Y8D8_inv pl=130n pw=800.0n nl=130n nw=800.0n
XI126 net186 VDDP VSS CENINT / S013LLLPSP_X256Y8D8_inv pl=130n pw=1.6u nl=130n nw=800.0n
XI127 CENINT VDDP VSS net186 / S013LLLPSP_X256Y8D8_inv pl=300n pw=250.00n nl=600n nw=250.00n
XI166 PRESACK1 VDDP VSS net273 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI129 net173 VDDP VSS net277 / S013LLLPSP_X256Y8D8_inv pl=130n pw=2u nl=130n nw=1.0u
XI130 net0334 VDDP VSS net281 / S013LLLPSP_X256Y8D8_inv pl=130n pw=4u nl=130n nw=2u
XI207 net277 VDDP VSS net0334 / S013LLLPSP_X256Y8D8_inv pl=130n pw=4u nl=130n nw=2u
XI133 FB_right VDDP VSS net285 / S013LLLPSP_X256Y8D8_inv pl=130n pw=1.6u nl=130n nw=1.6u
XI141 CLKLATCH VDDP VSS PRESACK1 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=20u nl=130.00n nw=10u
XI142 PRESACK1 VDDP VSS CLKLATCH / S013LLLPSP_X256Y8D8_inv pl=200.0n pw=250.00n nl=1u nw=250.00n
XI187 net0397 VDDP VSS SACK1_right / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=5u
XI144 net178 VDDP VSS ACTRCLK / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI145 ACTRCLK VDDP VSS ACTRCLKX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI146 net309 VDDP VSS DCTRCLKX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI147 net178 VDDP VSS net309 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=6u nl=130.00n nw=6u
XI148 net178 VDDP VSS DCTRCLK / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=10u nl=130.00n nw=5u
XI149 net0227 VDDP VSS net317 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI150 net317 VDDP VSS CLKD / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI152 net183 VDDP VSS SACK4 / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=5u
XI153 PRESACK1 VDDP VSS SACK1 / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=5u
XI156 PRESACK1 VDDP VSS INTCLKX / S013LLLPSP_X256Y8D8_inv pl=130n pw=10u nl=130n nw=10u
XI213 PRESACK1 VDDP VSS net0352 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
XI167 net273 VDDP VSS net337 / S013LLLPSP_X256Y8D8_inv pl=400n pw=800.0n nl=400n nw=800.0n
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_common_mode_Y8
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_common_mode_Y8 ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right DCTRCLK_right
+EMCLK FB_right FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0]
+FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] INTCLKX INTCLKX_right
+PXA[3] PXA[2] PXA[1] PXA[0] PXA_right[3] PXA_right[2] PXA_right[1] PXA_right[0] PXB[3] PXB[2]
+PXB[1] PXB[0] PXB_right[3] PXB_right[2] PXB_right[1] PXB_right[0] PXC[3] PXC[2] PXC[1] PXC[0]
+PXC_right[3] PXC_right[2] PXC_right[1] PXC_right[0] RDE S[1] S[0] SACK1 SACK1_right SACK4
+SACK4_right SM VDDP VMINE VSS WE WEN WE_right XA[8] XA[7]
+XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] XA[0] YA[2] YA[1] YA[0]
+YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] YX_right[7] YX_right[6]
+YX_right[5] YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0]
XICLKDRV ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX  DCTRCLKX_right DCTRCLK_right EMCLK FB_right INTCLKX INTCLKX_right S[1] S[0]  SACK1 SACK1_right SACK4 SACK4_right SM VDDP VMINE VSS WE WEN WE_right /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_CLKDRV_mode_V1
XI13 XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] XA[0] YA[2] YA[1] YA[0] CEN CLK  S[1] S[0] VDDP VSS WEN / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_ESDA14
XI19 XA[3] XA[4] ACTRCLK_right ACTRCLKX_right PXA_right[3] PXA_right[2]  PXA_right[1] PXA_right[0] RDE VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PXA
XPA XA[3] XA[4] ACTRCLK ACTRCLKX PXA[3] PXA[2] PXA[1] PXA[0] RDE VDDP VSS /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PXA
XI22 XA[7] XA[8] ACTRCLK_right ACTRCLKX_right PXC_right[3] PXC_right[2]  PXC_right[1] PXC_right[0] VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4
XI21 XA[5] XA[6] ACTRCLK_right ACTRCLKX_right PXB_right[3] PXB_right[2]  PXB_right[1] PXB_right[0] VDDP VSS / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4
XI10 XA[5] XA[6] ACTRCLK ACTRCLKX PXB[3] PXB[2] PXB[1] PXB[0] VDDP VSS /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4
XI11 XA[7] XA[8] ACTRCLK ACTRCLKX PXC[3] PXC[2] PXC[1] PXC[0] VDDP VSS /  S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_PX4
XI26 YA[0] YA[1] YA[2] ACTRCLK_right ACTRCLKX_right YX_right[7] YX_right[6]  YX_right[5] YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0] VDDP  VSS INTCLKX_right / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC
XI23 XA[0] XA[1] XA[2] ACTRCLK_right ACTRCLKX_right FCKX_right[7]  FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2]  FCKX_right[1] FCKX_right[0] VDDP VSS INTCLKX_right / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC
XI25 YA[0] YA[1] YA[2] ACTRCLK ACTRCLKX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]  YX[1] YX[0] VDDP VSS INTCLKX / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC
XIFPRE XA[0] XA[1] XA[2] ACTRCLK ACTRCLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4]  FCKX[3] FCKX[2] FCKX[1] FCKX[0] VDDP VSS INTCLKX / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FPREDEC
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11 FCKX PABC PABCX VDDP VSS WLL
MM1 WLL C VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS C / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=150.00n nw=1.5u
XI8 A VDDP VSS B / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=700.0n nl=130.00n nw=1u
XI114 A PABC PABCX VDDP VSS FCKX / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
MM0 WLL C VDDP VDDP P15LL W=2.5u L=150.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDDP VSS WLL[7] WLL[6] WLL[5] WLL[4] WLL[3] WLL[2] WLL[1]
+WLL[0]
XI156 PXA PXB PXC VDDP VSS net31 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLL[7] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLL[6] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLL[5] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLL[4] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLL[3] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLL[2] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLL[1] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLL[0] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_left_V0P11
XI111 net31 VDDP VSS PABC / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32left_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32left_V0P11 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXA_left[2]
+PXA_left[1] PXA_left[0] PXB_left[3] PXB_left[2] PXB_left[1] PXB_left[0] PXC_left[1] PXC_left[0] VDDP VSS
+WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248] WLL[247] WLL[246]
+WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238] WLL[237] WLL[236]
+WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226]
+WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217] WLL[216]
+WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208] WLL[207] WLL[206]
+WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198] WLL[197] WLL[196]
+WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186]
+WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177] WLL[176]
+WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168] WLL[167] WLL[166]
+WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158] WLL[157] WLL[156]
+WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146]
+WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137] WLL[136]
+WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128] WLL[127] WLL[126]
+WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118] WLL[117] WLL[116]
+WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106]
+WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97] WLL[96]
+WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88] WLL[87] WLL[86]
+WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78] WLL[77] WLL[76]
+WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66]
+WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57] WLL[56]
+WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48] WLL[47] WLL[46]
+WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38] WLL[37] WLL[36]
+WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26]
+WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17] WLL[16]
+WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8] WLL[7] WLL[6]
+WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0]
XIS013EELPSP_0 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[3]
+PXC_left[1] VDDP VSS WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249]
+WLL[248] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_1 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[3]
+PXC_left[1] VDDP VSS WLL[247] WLL[246] WLL[245] WLL[244] WLL[243] WLL[242] WLL[241]
+WLL[240] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_2 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[3]
+PXC_left[1] VDDP VSS WLL[239] WLL[238] WLL[237] WLL[236] WLL[235] WLL[234] WLL[233]
+WLL[232] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_3 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[3]
+PXC_left[1] VDDP VSS WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226] WLL[225]
+WLL[224] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_4 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[2]
+PXC_left[1] VDDP VSS WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217]
+WLL[216] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_5 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[2]
+PXC_left[1] VDDP VSS WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209]
+WLL[208] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_6 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[2]
+PXC_left[1] VDDP VSS WLL[207] WLL[206] WLL[205] WLL[204] WLL[203] WLL[202] WLL[201]
+WLL[200] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_7 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[2]
+PXC_left[1] VDDP VSS WLL[199] WLL[198] WLL[197] WLL[196] WLL[195] WLL[194] WLL[193]
+WLL[192] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_8 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[1]
+PXC_left[1] VDDP VSS WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186] WLL[185]
+WLL[184] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_9 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[1]
+PXC_left[1] VDDP VSS WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177]
+WLL[176] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_10 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[1]
+PXC_left[1] VDDP VSS WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169]
+WLL[168] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_11 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[1]
+PXC_left[1] VDDP VSS WLL[167] WLL[166] WLL[165] WLL[164] WLL[163] WLL[162] WLL[161]
+WLL[160] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_12 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[0]
+PXC_left[1] VDDP VSS WLL[159] WLL[158] WLL[157] WLL[156] WLL[155] WLL[154] WLL[153]
+WLL[152] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_13 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[0]
+PXC_left[1] VDDP VSS WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146] WLL[145]
+WLL[144] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_14 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[0]
+PXC_left[1] VDDP VSS WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137]
+WLL[136] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_15 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[0]
+PXC_left[1] VDDP VSS WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129]
+WLL[128] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_16 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[3]
+PXC_left[0] VDDP VSS WLL[127] WLL[126] WLL[125] WLL[124] WLL[123] WLL[122] WLL[121]
+WLL[120] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_17 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[3]
+PXC_left[0] VDDP VSS WLL[119] WLL[118] WLL[117] WLL[116] WLL[115] WLL[114] WLL[113]
+WLL[112] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_18 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[3]
+PXC_left[0] VDDP VSS WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106] WLL[105]
+WLL[104] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_19 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[3]
+PXC_left[0] VDDP VSS WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97]
+WLL[96] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_20 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[2]
+PXC_left[0] VDDP VSS WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89]
+WLL[88] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_21 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[2]
+PXC_left[0] VDDP VSS WLL[87] WLL[86] WLL[85] WLL[84] WLL[83] WLL[82] WLL[81]
+WLL[80] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_22 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[2]
+PXC_left[0] VDDP VSS WLL[79] WLL[78] WLL[77] WLL[76] WLL[75] WLL[74] WLL[73]
+WLL[72] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_23 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[2]
+PXC_left[0] VDDP VSS WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66] WLL[65]
+WLL[64] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_24 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[1]
+PXC_left[0] VDDP VSS WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57]
+WLL[56] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_25 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[1]
+PXC_left[0] VDDP VSS WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49]
+WLL[48] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_26 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[1]
+PXC_left[0] VDDP VSS WLL[47] WLL[46] WLL[45] WLL[44] WLL[43] WLL[42] WLL[41]
+WLL[40] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_27 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[1]
+PXC_left[0] VDDP VSS WLL[39] WLL[38] WLL[37] WLL[36] WLL[35] WLL[34] WLL[33]
+WLL[32] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_28 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[3] PXB_left[0]
+PXC_left[0] VDDP VSS WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26] WLL[25]
+WLL[24] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_29 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[2] PXB_left[0]
+PXC_left[0] VDDP VSS WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17]
+WLL[16] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_30 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[1] PXB_left[0]
+PXC_left[0] VDDP VSS WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9]
+WLL[8] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
XIS013EELPSP_31 FCKX_left[7] FCKX_left[6] FCKX_left[5] FCKX_left[4] FCKX_left[3] FCKX_left[2] FCKX_left[1] FCKX_left[0] PXA_left[0] PXB_left[0]
+PXC_left[0] VDDP VSS WLL[7] WLL[6] WLL[5] WLL[4] WLL[3] WLL[2] WLL[1]
+WLL[0] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_left_V0P11
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11 FCKX PABC PABCX VDDP VSS WLR
MM2 WLR net46 VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS net46 / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=150.00n nw=1.5u
XI8 A VDDP VSS B / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=700.0n nl=130.00n nw=1u
XI114 A PABC PABCX VDDP VSS FCKX / S013LLLPSP_X256Y8D8_tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
MM3 WLR net46 VDDP VDDP P15LL W=2.5u L=150.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDDP VSS WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1]
+WLR[0]
XI156 PXA PXB PXC VDDP VSS net31 / S013LLLPSP_X256Y8D8_nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLR[7] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLR[6] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLR[5] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLR[4] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLR[3] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLR[2] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLR[1] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLR[0] / S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_FDEC_right_V0P11
XI111 net31 VDDP VSS PABC / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / S013LLLPSP_X256Y8D8_inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32right_V0P11
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32right_V0P11 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXA_right[2]
+PXA_right[1] PXA_right[0] PXB_right[3] PXB_right[2] PXB_right[1] PXB_right[0] PXC_right[1] PXC_right[0] VDDP VSS
+WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250] WLR[249] WLR[248] WLR[247] WLR[246]
+WLR[245] WLR[244] WLR[243] WLR[242] WLR[241] WLR[240] WLR[239] WLR[238] WLR[237] WLR[236]
+WLR[235] WLR[234] WLR[233] WLR[232] WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226]
+WLR[225] WLR[224] WLR[223] WLR[222] WLR[221] WLR[220] WLR[219] WLR[218] WLR[217] WLR[216]
+WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210] WLR[209] WLR[208] WLR[207] WLR[206]
+WLR[205] WLR[204] WLR[203] WLR[202] WLR[201] WLR[200] WLR[199] WLR[198] WLR[197] WLR[196]
+WLR[195] WLR[194] WLR[193] WLR[192] WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186]
+WLR[185] WLR[184] WLR[183] WLR[182] WLR[181] WLR[180] WLR[179] WLR[178] WLR[177] WLR[176]
+WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170] WLR[169] WLR[168] WLR[167] WLR[166]
+WLR[165] WLR[164] WLR[163] WLR[162] WLR[161] WLR[160] WLR[159] WLR[158] WLR[157] WLR[156]
+WLR[155] WLR[154] WLR[153] WLR[152] WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146]
+WLR[145] WLR[144] WLR[143] WLR[142] WLR[141] WLR[140] WLR[139] WLR[138] WLR[137] WLR[136]
+WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130] WLR[129] WLR[128] WLR[127] WLR[126]
+WLR[125] WLR[124] WLR[123] WLR[122] WLR[121] WLR[120] WLR[119] WLR[118] WLR[117] WLR[116]
+WLR[115] WLR[114] WLR[113] WLR[112] WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106]
+WLR[105] WLR[104] WLR[103] WLR[102] WLR[101] WLR[100] WLR[99] WLR[98] WLR[97] WLR[96]
+WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90] WLR[89] WLR[88] WLR[87] WLR[86]
+WLR[85] WLR[84] WLR[83] WLR[82] WLR[81] WLR[80] WLR[79] WLR[78] WLR[77] WLR[76]
+WLR[75] WLR[74] WLR[73] WLR[72] WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66]
+WLR[65] WLR[64] WLR[63] WLR[62] WLR[61] WLR[60] WLR[59] WLR[58] WLR[57] WLR[56]
+WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50] WLR[49] WLR[48] WLR[47] WLR[46]
+WLR[45] WLR[44] WLR[43] WLR[42] WLR[41] WLR[40] WLR[39] WLR[38] WLR[37] WLR[36]
+WLR[35] WLR[34] WLR[33] WLR[32] WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26]
+WLR[25] WLR[24] WLR[23] WLR[22] WLR[21] WLR[20] WLR[19] WLR[18] WLR[17] WLR[16]
+WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10] WLR[9] WLR[8] WLR[7] WLR[6]
+WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0]
XIS013EELPSP_0 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[3]
+PXC_right[1] VDDP VSS WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250] WLR[249]
+WLR[248] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_1 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[3]
+PXC_right[1] VDDP VSS WLR[247] WLR[246] WLR[245] WLR[244] WLR[243] WLR[242] WLR[241]
+WLR[240] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_2 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[3]
+PXC_right[1] VDDP VSS WLR[239] WLR[238] WLR[237] WLR[236] WLR[235] WLR[234] WLR[233]
+WLR[232] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_3 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[3]
+PXC_right[1] VDDP VSS WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226] WLR[225]
+WLR[224] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_4 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[2]
+PXC_right[1] VDDP VSS WLR[223] WLR[222] WLR[221] WLR[220] WLR[219] WLR[218] WLR[217]
+WLR[216] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_5 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[2]
+PXC_right[1] VDDP VSS WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210] WLR[209]
+WLR[208] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_6 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[2]
+PXC_right[1] VDDP VSS WLR[207] WLR[206] WLR[205] WLR[204] WLR[203] WLR[202] WLR[201]
+WLR[200] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_7 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[2]
+PXC_right[1] VDDP VSS WLR[199] WLR[198] WLR[197] WLR[196] WLR[195] WLR[194] WLR[193]
+WLR[192] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_8 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[1]
+PXC_right[1] VDDP VSS WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186] WLR[185]
+WLR[184] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_9 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[1]
+PXC_right[1] VDDP VSS WLR[183] WLR[182] WLR[181] WLR[180] WLR[179] WLR[178] WLR[177]
+WLR[176] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_10 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[1]
+PXC_right[1] VDDP VSS WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170] WLR[169]
+WLR[168] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_11 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[1]
+PXC_right[1] VDDP VSS WLR[167] WLR[166] WLR[165] WLR[164] WLR[163] WLR[162] WLR[161]
+WLR[160] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_12 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[0]
+PXC_right[1] VDDP VSS WLR[159] WLR[158] WLR[157] WLR[156] WLR[155] WLR[154] WLR[153]
+WLR[152] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_13 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[0]
+PXC_right[1] VDDP VSS WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146] WLR[145]
+WLR[144] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_14 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[0]
+PXC_right[1] VDDP VSS WLR[143] WLR[142] WLR[141] WLR[140] WLR[139] WLR[138] WLR[137]
+WLR[136] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_15 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[0]
+PXC_right[1] VDDP VSS WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130] WLR[129]
+WLR[128] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_16 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[3]
+PXC_right[0] VDDP VSS WLR[127] WLR[126] WLR[125] WLR[124] WLR[123] WLR[122] WLR[121]
+WLR[120] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_17 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[3]
+PXC_right[0] VDDP VSS WLR[119] WLR[118] WLR[117] WLR[116] WLR[115] WLR[114] WLR[113]
+WLR[112] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_18 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[3]
+PXC_right[0] VDDP VSS WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106] WLR[105]
+WLR[104] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_19 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[3]
+PXC_right[0] VDDP VSS WLR[103] WLR[102] WLR[101] WLR[100] WLR[99] WLR[98] WLR[97]
+WLR[96] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_20 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[2]
+PXC_right[0] VDDP VSS WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90] WLR[89]
+WLR[88] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_21 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[2]
+PXC_right[0] VDDP VSS WLR[87] WLR[86] WLR[85] WLR[84] WLR[83] WLR[82] WLR[81]
+WLR[80] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_22 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[2]
+PXC_right[0] VDDP VSS WLR[79] WLR[78] WLR[77] WLR[76] WLR[75] WLR[74] WLR[73]
+WLR[72] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_23 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[2]
+PXC_right[0] VDDP VSS WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66] WLR[65]
+WLR[64] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_24 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[1]
+PXC_right[0] VDDP VSS WLR[63] WLR[62] WLR[61] WLR[60] WLR[59] WLR[58] WLR[57]
+WLR[56] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_25 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[1]
+PXC_right[0] VDDP VSS WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50] WLR[49]
+WLR[48] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_26 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[1]
+PXC_right[0] VDDP VSS WLR[47] WLR[46] WLR[45] WLR[44] WLR[43] WLR[42] WLR[41]
+WLR[40] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_27 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[1]
+PXC_right[0] VDDP VSS WLR[39] WLR[38] WLR[37] WLR[36] WLR[35] WLR[34] WLR[33]
+WLR[32] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_28 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXB_right[0]
+PXC_right[0] VDDP VSS WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26] WLR[25]
+WLR[24] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_29 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[2] PXB_right[0]
+PXC_right[0] VDDP VSS WLR[23] WLR[22] WLR[21] WLR[20] WLR[19] WLR[18] WLR[17]
+WLR[16] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_30 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[1] PXB_right[0]
+PXC_right[0] VDDP VSS WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10] WLR[9]
+WLR[8] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
XIS013EELPSP_31 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[0] PXB_right[0]
+PXC_right[0] VDDP VSS WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1]
+WLR[0] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_XDEC_right_V0P11
.ENDS

************************************************************************
* Library Name: SMIC_MEMORY
* Cell Name:    S013LLLPSP_X256Y8D8
* View Name:    schematic
************************************************************************

.SUBCKT S013LLLPSP_X256Y8D8 WEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] D[7]
+D[6] D[5] D[4] D[3] D[2] D[1] D[0] CLK CEN A[10]
+A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+VDDP VDDC VSS
XIS013EELPSP_0 TIEH VDDP VSS S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieH
XIS013EELPSP_1 TIEL VDDP VSS S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_TieL
XIS013EELPSP_2 TIEL TIEL TIEL TIEL D[7] D[6] D[5] D[4] DBL_right DCTRCLK_right
+DCTRCLKX_right Q[7] Q[6] Q[5] Q[4] RWLR VSS SACK1_right SACK4_right STWL_right
+VDDP VDDC VSS WE_right WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250]
+WLR[249] WLR[248] WLR[247] WLR[246] WLR[245] WLR[244] WLR[243] WLR[242] WLR[241] WLR[240]
+WLR[239] WLR[238] WLR[237] WLR[236] WLR[235] WLR[234] WLR[233] WLR[232] WLR[231] WLR[230]
+WLR[229] WLR[228] WLR[227] WLR[226] WLR[225] WLR[224] WLR[223] WLR[222] WLR[221] WLR[220]
+WLR[219] WLR[218] WLR[217] WLR[216] WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210]
+WLR[209] WLR[208] WLR[207] WLR[206] WLR[205] WLR[204] WLR[203] WLR[202] WLR[201] WLR[200]
+WLR[199] WLR[198] WLR[197] WLR[196] WLR[195] WLR[194] WLR[193] WLR[192] WLR[191] WLR[190]
+WLR[189] WLR[188] WLR[187] WLR[186] WLR[185] WLR[184] WLR[183] WLR[182] WLR[181] WLR[180]
+WLR[179] WLR[178] WLR[177] WLR[176] WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170]
+WLR[169] WLR[168] WLR[167] WLR[166] WLR[165] WLR[164] WLR[163] WLR[162] WLR[161] WLR[160]
+WLR[159] WLR[158] WLR[157] WLR[156] WLR[155] WLR[154] WLR[153] WLR[152] WLR[151] WLR[150]
+WLR[149] WLR[148] WLR[147] WLR[146] WLR[145] WLR[144] WLR[143] WLR[142] WLR[141] WLR[140]
+WLR[139] WLR[138] WLR[137] WLR[136] WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130]
+WLR[129] WLR[128] WLR[127] WLR[126] WLR[125] WLR[124] WLR[123] WLR[122] WLR[121] WLR[120]
+WLR[119] WLR[118] WLR[117] WLR[116] WLR[115] WLR[114] WLR[113] WLR[112] WLR[111] WLR[110]
+WLR[109] WLR[108] WLR[107] WLR[106] WLR[105] WLR[104] WLR[103] WLR[102] WLR[101] WLR[100]
+WLR[99] WLR[98] WLR[97] WLR[96] WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90]
+WLR[89] WLR[88] WLR[87] WLR[86] WLR[85] WLR[84] WLR[83] WLR[82] WLR[81] WLR[80]
+WLR[79] WLR[78] WLR[77] WLR[76] WLR[75] WLR[74] WLR[73] WLR[72] WLR[71] WLR[70]
+WLR[69] WLR[68] WLR[67] WLR[66] WLR[65] WLR[64] WLR[63] WLR[62] WLR[61] WLR[60]
+WLR[59] WLR[58] WLR[57] WLR[56] WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50]
+WLR[49] WLR[48] WLR[47] WLR[46] WLR[45] WLR[44] WLR[43] WLR[42] WLR[41] WLR[40]
+WLR[39] WLR[38] WLR[37] WLR[36] WLR[35] WLR[34] WLR[33] WLR[32] WLR[31] WLR[30]
+WLR[29] WLR[28] WLR[27] WLR[26] WLR[25] WLR[24] WLR[23] WLR[22] WLR[21] WLR[20]
+WLR[19] WLR[18] WLR[17] WLR[16] WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10]
+WLR[9] WLR[8] WLR[7] WLR[6] WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0]
+YX_right[7] YX_right[6] YX_right[5] YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_right
XIS013EELPSP_3 TIEL TIEL TIEL TIEL D[3] D[2] D[1] D[0] DCTRCLK DCTRCLKX
+Q[3] Q[2] Q[1] Q[0] RWLL VSS SACK1 SACK4 VDDP VDDC
+VSS WE WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248]
+WLL[247] WLL[246] WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238]
+WLL[237] WLL[236] WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228]
+WLL[227] WLL[226] WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218]
+WLL[217] WLL[216] WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208]
+WLL[207] WLL[206] WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198]
+WLL[197] WLL[196] WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188]
+WLL[187] WLL[186] WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178]
+WLL[177] WLL[176] WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168]
+WLL[167] WLL[166] WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158]
+WLL[157] WLL[156] WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148]
+WLL[147] WLL[146] WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138]
+WLL[137] WLL[136] WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128]
+WLL[127] WLL[126] WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118]
+WLL[117] WLL[116] WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108]
+WLL[107] WLL[106] WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98]
+WLL[97] WLL[96] WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88]
+WLL[87] WLL[86] WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78]
+WLL[77] WLL[76] WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68]
+WLL[67] WLL[66] WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58]
+WLL[57] WLL[56] WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48]
+WLL[47] WLL[46] WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38]
+WLL[37] WLL[36] WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28]
+WLL[27] WLL[26] WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18]
+WLL[17] WLL[16] WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8]
+WLL[7] WLL[6] WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0] YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] S013LLLPSP_X256Y8D8_S013EELPSP_array_X256Y8D4BWEN_left
XIS013EELPSP_4 ACTRCLK ACTRCLKX TIEL RWLL VDDP VSS INTCLKX S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_left
XIS013EELPSP_5 ACTRCLK_right ACTRCLKX_right TIEL RWLR VDDP VSS INTCLKX_right S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_RWL_DEC_right
XIS013EELPSP_6 DBL_right EMCLK STWL_right VDDP VSS S013LLLPSP_X256Y8D8_S013EELPSP_SOP01
XIS013EELPSP_7 ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right DCTRCLK_right
+EMCLK DBL_right FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0]
+FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] INTCLKX INTCLKX_right
+PXA[3] PXA[2] PXA[1] PXA[0] PXA_right[3] PXA_right[2] PXA_right[1] PXA_right[0] PXB[3] PXB[2]
+PXB[1] PXB[0] PXB_right[3] PXB_right[2] PXB_right[1] PXB_right[0] PXC[3] PXC[2] PXC[1] PXC[0]
+PXC_right[3] PXC_right[2] PXC_right[1] PXC_right[0] TIEL TIEH TIEH SACK1 SACK1_right SACK4
+SACK4_right TIEL VDDP TIEL VSS WE WEN WE_right TIEL A[10]
+A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+YX[7] YX[6] YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] YX_right[7] YX_right[6]
+YX_right[5] YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0] S013LLLPSP_X256Y8D8_S013EELPSP_LEAFCELL_Logic_common_mode_Y8
XIS013EELPSP_8 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2]
+PXA[1] PXA[0] PXB[3] PXB[2] PXB[1] PXB[0] PXC[1] PXC[0] VDDP VSS
+WLL[255] WLL[254] WLL[253] WLL[252] WLL[251] WLL[250] WLL[249] WLL[248] WLL[247] WLL[246]
+WLL[245] WLL[244] WLL[243] WLL[242] WLL[241] WLL[240] WLL[239] WLL[238] WLL[237] WLL[236]
+WLL[235] WLL[234] WLL[233] WLL[232] WLL[231] WLL[230] WLL[229] WLL[228] WLL[227] WLL[226]
+WLL[225] WLL[224] WLL[223] WLL[222] WLL[221] WLL[220] WLL[219] WLL[218] WLL[217] WLL[216]
+WLL[215] WLL[214] WLL[213] WLL[212] WLL[211] WLL[210] WLL[209] WLL[208] WLL[207] WLL[206]
+WLL[205] WLL[204] WLL[203] WLL[202] WLL[201] WLL[200] WLL[199] WLL[198] WLL[197] WLL[196]
+WLL[195] WLL[194] WLL[193] WLL[192] WLL[191] WLL[190] WLL[189] WLL[188] WLL[187] WLL[186]
+WLL[185] WLL[184] WLL[183] WLL[182] WLL[181] WLL[180] WLL[179] WLL[178] WLL[177] WLL[176]
+WLL[175] WLL[174] WLL[173] WLL[172] WLL[171] WLL[170] WLL[169] WLL[168] WLL[167] WLL[166]
+WLL[165] WLL[164] WLL[163] WLL[162] WLL[161] WLL[160] WLL[159] WLL[158] WLL[157] WLL[156]
+WLL[155] WLL[154] WLL[153] WLL[152] WLL[151] WLL[150] WLL[149] WLL[148] WLL[147] WLL[146]
+WLL[145] WLL[144] WLL[143] WLL[142] WLL[141] WLL[140] WLL[139] WLL[138] WLL[137] WLL[136]
+WLL[135] WLL[134] WLL[133] WLL[132] WLL[131] WLL[130] WLL[129] WLL[128] WLL[127] WLL[126]
+WLL[125] WLL[124] WLL[123] WLL[122] WLL[121] WLL[120] WLL[119] WLL[118] WLL[117] WLL[116]
+WLL[115] WLL[114] WLL[113] WLL[112] WLL[111] WLL[110] WLL[109] WLL[108] WLL[107] WLL[106]
+WLL[105] WLL[104] WLL[103] WLL[102] WLL[101] WLL[100] WLL[99] WLL[98] WLL[97] WLL[96]
+WLL[95] WLL[94] WLL[93] WLL[92] WLL[91] WLL[90] WLL[89] WLL[88] WLL[87] WLL[86]
+WLL[85] WLL[84] WLL[83] WLL[82] WLL[81] WLL[80] WLL[79] WLL[78] WLL[77] WLL[76]
+WLL[75] WLL[74] WLL[73] WLL[72] WLL[71] WLL[70] WLL[69] WLL[68] WLL[67] WLL[66]
+WLL[65] WLL[64] WLL[63] WLL[62] WLL[61] WLL[60] WLL[59] WLL[58] WLL[57] WLL[56]
+WLL[55] WLL[54] WLL[53] WLL[52] WLL[51] WLL[50] WLL[49] WLL[48] WLL[47] WLL[46]
+WLL[45] WLL[44] WLL[43] WLL[42] WLL[41] WLL[40] WLL[39] WLL[38] WLL[37] WLL[36]
+WLL[35] WLL[34] WLL[33] WLL[32] WLL[31] WLL[30] WLL[29] WLL[28] WLL[27] WLL[26]
+WLL[25] WLL[24] WLL[23] WLL[22] WLL[21] WLL[20] WLL[19] WLL[18] WLL[17] WLL[16]
+WLL[15] WLL[14] WLL[13] WLL[12] WLL[11] WLL[10] WLL[9] WLL[8] WLL[7] WLL[6]
+WLL[5] WLL[4] WLL[3] WLL[2] WLL[1] WLL[0] S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32left_V0P11
XIS013EELPSP_9 FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] PXA_right[3] PXA_right[2]
+PXA_right[1] PXA_right[0] PXB_right[3] PXB_right[2] PXB_right[1] PXB_right[0] PXC_right[1] PXC_right[0] VDDP VSS
+WLR[255] WLR[254] WLR[253] WLR[252] WLR[251] WLR[250] WLR[249] WLR[248] WLR[247] WLR[246]
+WLR[245] WLR[244] WLR[243] WLR[242] WLR[241] WLR[240] WLR[239] WLR[238] WLR[237] WLR[236]
+WLR[235] WLR[234] WLR[233] WLR[232] WLR[231] WLR[230] WLR[229] WLR[228] WLR[227] WLR[226]
+WLR[225] WLR[224] WLR[223] WLR[222] WLR[221] WLR[220] WLR[219] WLR[218] WLR[217] WLR[216]
+WLR[215] WLR[214] WLR[213] WLR[212] WLR[211] WLR[210] WLR[209] WLR[208] WLR[207] WLR[206]
+WLR[205] WLR[204] WLR[203] WLR[202] WLR[201] WLR[200] WLR[199] WLR[198] WLR[197] WLR[196]
+WLR[195] WLR[194] WLR[193] WLR[192] WLR[191] WLR[190] WLR[189] WLR[188] WLR[187] WLR[186]
+WLR[185] WLR[184] WLR[183] WLR[182] WLR[181] WLR[180] WLR[179] WLR[178] WLR[177] WLR[176]
+WLR[175] WLR[174] WLR[173] WLR[172] WLR[171] WLR[170] WLR[169] WLR[168] WLR[167] WLR[166]
+WLR[165] WLR[164] WLR[163] WLR[162] WLR[161] WLR[160] WLR[159] WLR[158] WLR[157] WLR[156]
+WLR[155] WLR[154] WLR[153] WLR[152] WLR[151] WLR[150] WLR[149] WLR[148] WLR[147] WLR[146]
+WLR[145] WLR[144] WLR[143] WLR[142] WLR[141] WLR[140] WLR[139] WLR[138] WLR[137] WLR[136]
+WLR[135] WLR[134] WLR[133] WLR[132] WLR[131] WLR[130] WLR[129] WLR[128] WLR[127] WLR[126]
+WLR[125] WLR[124] WLR[123] WLR[122] WLR[121] WLR[120] WLR[119] WLR[118] WLR[117] WLR[116]
+WLR[115] WLR[114] WLR[113] WLR[112] WLR[111] WLR[110] WLR[109] WLR[108] WLR[107] WLR[106]
+WLR[105] WLR[104] WLR[103] WLR[102] WLR[101] WLR[100] WLR[99] WLR[98] WLR[97] WLR[96]
+WLR[95] WLR[94] WLR[93] WLR[92] WLR[91] WLR[90] WLR[89] WLR[88] WLR[87] WLR[86]
+WLR[85] WLR[84] WLR[83] WLR[82] WLR[81] WLR[80] WLR[79] WLR[78] WLR[77] WLR[76]
+WLR[75] WLR[74] WLR[73] WLR[72] WLR[71] WLR[70] WLR[69] WLR[68] WLR[67] WLR[66]
+WLR[65] WLR[64] WLR[63] WLR[62] WLR[61] WLR[60] WLR[59] WLR[58] WLR[57] WLR[56]
+WLR[55] WLR[54] WLR[53] WLR[52] WLR[51] WLR[50] WLR[49] WLR[48] WLR[47] WLR[46]
+WLR[45] WLR[44] WLR[43] WLR[42] WLR[41] WLR[40] WLR[39] WLR[38] WLR[37] WLR[36]
+WLR[35] WLR[34] WLR[33] WLR[32] WLR[31] WLR[30] WLR[29] WLR[28] WLR[27] WLR[26]
+WLR[25] WLR[24] WLR[23] WLR[22] WLR[21] WLR[20] WLR[19] WLR[18] WLR[17] WLR[16]
+WLR[15] WLR[14] WLR[13] WLR[12] WLR[11] WLR[10] WLR[9] WLR[8] WLR[7] WLR[6]
+WLR[5] WLR[4] WLR[3] WLR[2] WLR[1] WLR[0] S013LLLPSP_X256Y8D8_S013EELPSP_XDEC32right_V0P11
.ENDS
