# Copyright (c) 2024 SMIC
# Filename   : S013LLLPSP_X256Y8D8.lef
# IP code    : S013LLLPSP
# Version    : v0p2
# CreateDate : Sep 19, 2024

# Name: Single-Port Low Power SRAM, SMIC 0.13um  EE Process
# Configuration: -instname S013LLLPSP_X256Y8D8 -rows 256 -bits 8 -mux 8 
# Redundancy: Off
# Bit-Write: Off

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO S013LLLPSP_X256Y8D8
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 182.34 BY 559.045 ;
 PIN Q[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 3.965 0 4.165 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[0]
 PIN D[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 5.555 0 5.755 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[0]
 PIN D[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 20.745 0 20.945 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[1]
 PIN Q[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 22.335 0 22.535 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[1]
 PIN Q[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 26.305 0 26.505 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[2]
 PIN D[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 27.895 0 28.095 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[2]
 PIN D[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 43.085 0 43.285 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[3]
 PIN Q[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 44.675 0 44.875 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[3]
 PIN WEN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 57.37 0 57.57 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END WEN
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 79.3 0 79.55 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END CLK
 PIN CEN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 80.885 0 81.135 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END CEN
 PIN A[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 96.22 0 96.42 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[7]
 PIN A[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 98.535 0 98.735 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[6]
 PIN A[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 101.77 0 101.97 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[9]
 PIN A[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 104.085 0 104.285 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[8]
 PIN A[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 109.635 0 109.835 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[10]
 PIN A[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 114.2 0 114.4 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[3]
 PIN A[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 116.44 0 116.64 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[5]
 PIN A[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 119.8 0 120 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[4]
 PIN A[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 124.21 0 124.41 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[0]
 PIN A[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 125.33 0 125.53 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[2]
 PIN A[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 127.61 0 127.81 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END A[1]
 PIN Q[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 137.465 0 137.665 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[4]
 PIN D[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 139.055 0 139.255 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[4]
 PIN D[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 154.245 0 154.445 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[5]
 PIN Q[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 155.835 0 156.035 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[5]
 PIN Q[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 159.805 0 160.005 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[6]
 PIN D[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 161.395 0 161.595 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[6]
 PIN D[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 176.585 0 176.785 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END D[7]
 PIN Q[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M2 ;
 RECT 178.175 0 178.375 0.5 ;
 END
 ANTENNAGATEAREA 0.208 ;
 ANTENNADIFFAREA 0.1736 ;
 END Q[7]
 PIN VDDP
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 52.44 0 53.04 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 57.045 0 57.645 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 60.645 0 61.245 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 64.245 0 64.845 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 67.845 0 68.445 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 71.445 0 72.045 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 75.045 0 75.645 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 78.645 0 79.245 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 82.245 0 82.845 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 85.845 0 86.445 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 89.445 0 90.045 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 92.295 0 92.895 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 95.895 0 96.495 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 99.495 0 100.095 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 103.095 0 103.695 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 106.695 0 107.295 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 110.295 0 110.895 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 113.895 0 114.495 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 117.495 0 118.095 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 121.095 0 121.695 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 124.695 0 125.295 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 129.3 0 129.9 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 0.635 0 1.235 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 2.925 0 3.525 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 12.335 0 12.935 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 13.565 0 14.165 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 22.975 0 23.575 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 25.265 0 25.865 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 34.675 0 35.275 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 35.905 0 36.505 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 45.315 0 45.915 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 47.605 0 48.205 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 134.135 0 134.735 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 136.425 0 137.025 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 145.835 0 146.435 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 147.065 0 147.665 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 156.475 0 157.075 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 158.765 0 159.365 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 168.175 0 168.775 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 169.405 0 170.005 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 178.815 0 179.415 559.045 ; 
 END 
 PORT
 LAYER M4 ;
 RECT 181.105 0 181.705 559.045 ; 
 END 
 END VDDP
 PIN VDDC
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 7.015 0 7.615 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 8.245 0 8.845 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 17.655 0 18.255 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 18.885 0 19.485 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 29.355 0 29.955 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 30.585 0 31.185 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 39.995 0 40.595 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 41.225 0 41.825 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 140.515 0 141.115 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 141.745 0 142.345 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 151.155 0 151.755 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 152.385 0 152.985 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 162.855 0 163.455 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 164.085 0 164.685 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 173.495 0 174.095 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 174.725 0 175.325 559.045 ;    
 END 
 END VDDC
 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 55.195 0 55.795 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 58.845 0 59.445 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 62.445 0 63.045 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 66.045 0 66.645 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 69.645 0 70.245 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 73.245 0 73.845 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 76.845 0 77.445 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 80.445 0 81.045 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 84.045 0 84.645 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 87.645 0 88.245 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 94.095 0 94.695 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 97.695 0 98.295 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 101.295 0 101.895 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 104.895 0 105.495 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 108.495 0 109.095 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 112.095 0 112.695 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 115.695 0 116.295 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 119.295 0 119.895 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 122.895 0 123.495 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 126.545 0 127.145 559.045 ;      
 END
 PORT
 LAYER M4 ;
 RECT 1.78 0 2.38 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 4.355 0 4.955 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 5.585 0 6.185 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 9.675 0 10.275 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.905 0 11.505 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 14.995 0 15.595 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 16.225 0 16.825 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 20.315 0 20.915 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 21.545 0 22.145 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 24.12 0 24.72 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 26.695 0 27.295 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 27.925 0 28.525 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 32.015 0 32.615 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 33.245 0 33.845 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 37.335 0 37.935 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 38.565 0 39.165 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 42.655 0 43.255 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 43.885 0 44.485 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 46.46 0 47.06 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 135.28 0 135.88 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 137.855 0 138.455 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 139.085 0 139.685 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 143.175 0 143.775 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 144.405 0 145.005 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 148.495 0 149.095 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 149.725 0 150.325 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 153.815 0 154.415 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 155.045 0 155.645 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 157.62 0 158.22 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 160.195 0 160.795 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 161.425 0 162.025 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 165.515 0 166.115 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 166.745 0 167.345 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 170.835 0 171.435 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 172.065 0 172.665 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 176.155 0 176.755 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 177.385 0 177.985 559.045 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 179.96 0 180.56 559.045 ;    
 END 
 END VSS
 OBS
 LAYER M2 ;
 RECT 0 0 3.765 0.7 ;
 RECT 4.365 0 5.355 0.7 ;
 RECT 5.955 0 20.545 0.7 ;
 RECT 21.145 0 22.135 0.7 ;
 RECT 22.735 0 26.105 0.7 ;
 RECT 26.705 0 27.695 0.7 ;
 RECT 28.295 0 42.885 0.7 ;
 RECT 43.485 0 44.475 0.7 ;
 RECT 45.075 0 57.17 0.7 ;
 RECT 57.77 0 79.1 0.7 ;
 RECT 79.75 0 80.685 0.7 ;
 RECT 81.335 0 96.02 0.7 ;
 RECT 96.62 0 98.335 0.7 ;
 RECT 98.935 0 101.57 0.7 ;
 RECT 102.17 0 103.885 0.7 ;
 RECT 104.485 0 109.435 0.7 ;
 RECT 110.035 0 114 0.7 ;
 RECT 114.6 0 116.24 0.7 ;
 RECT 116.84 0 119.6 0.7 ;
 RECT 120.2 0 124.01 0.7 ;
 RECT 124.61 0 125.13 0.7 ;
 RECT 125.73 0 127.41 0.7 ;
 RECT 128.01 0 137.265 0.7 ;
 RECT 137.865 0 138.855 0.7 ;
 RECT 139.455 0 154.045 0.7 ;
 RECT 154.645 0 155.635 0.7 ;
 RECT 156.235 0 159.605 0.7 ;
 RECT 160.205 0 161.195 0.7 ;
 RECT 161.795 0 176.385 0.7 ;
 RECT 176.985 0 177.975 0.7 ;
 RECT  178.575 0 182.34 0.7 ;
 RECT  0 559.045 182.34 558.345 ;
 RECT 0 0.7 182.34 558.345 ;
 LAYER M1 ;
 RECT 0 0 182.34 559.045 ;
 LAYER M3 ;
 RECT 0 0 182.34 559.045 ;
 LAYER M4 ;
 RECT 0 0 0.385 559.045 ;
 RECT 3.775 0 4.105 559.045 ;
 RECT 6.435 0 6.765 559.045 ;
 RECT 9.095 0 9.425 559.045 ;
 RECT 11.755 0 12.085 559.045 ;
 RECT 14.415 0 14.745 559.045 ;
 RECT 17.075 0 17.405 559.045 ;
 RECT 19.735 0 20.065 559.045 ;
 RECT 22.395 0 22.725 559.045 ;
 RECT 26.115 0 26.445 559.045 ;
 RECT 28.775 0 29.105 559.045 ;
 RECT 31.435 0 31.765 559.045 ;
 RECT 34.095 0 34.425 559.045 ;
 RECT 36.755 0 37.085 559.045 ;
 RECT 39.415 0 39.745 559.045 ;
 RECT 42.075 0 42.405 559.045 ;
 RECT 44.735 0 45.065 559.045 ;
 RECT 48.455 0 52.19 559.045 ;
 RECT 53.29 0 54.945 559.045 ;
 RECT 56.045 0 56.795 559.045 ;
 RECT 57.895 0 58.595 559.045 ;
 RECT 59.695 0 60.395 559.045 ;
 RECT 61.495 0 62.195 559.045 ;
 RECT 63.295 0 63.995 559.045 ;
 RECT 65.095 0 65.795 559.045 ;
 RECT 66.895 0 67.595 559.045 ;
 RECT 68.695 0 69.395 559.045 ;
 RECT 70.495 0 71.195 559.045 ;
 RECT 72.295 0 72.995 559.045 ;
 RECT 74.095 0 74.795 559.045 ;
 RECT 75.895 0 76.595 559.045 ;
 RECT 77.695 0 78.395 559.045 ;
 RECT 79.495 0 80.195 559.045 ;
 RECT 81.295 0 81.995 559.045 ;
 RECT 83.095 0 83.795 559.045 ;
 RECT 84.895 0 85.595 559.045 ;
 RECT 86.695 0 87.395 559.045 ;
 RECT 88.495 0 89.195 559.045 ;
 RECT 90.295 0 92.045 559.045 ;
 RECT 93.145 0 93.845 559.045 ;
 RECT 94.945 0 95.645 559.045 ;
 RECT 96.745 0 97.445 559.045 ;
 RECT 98.545 0 99.245 559.045 ;
 RECT 100.345 0 101.045 559.045 ;
 RECT 102.145 0 102.845 559.045 ;
 RECT 103.945 0 104.645 559.045 ;
 RECT 105.745 0 106.445 559.045 ;
 RECT 107.545 0 108.245 559.045 ;
 RECT 109.345 0 110.045 559.045 ;
 RECT 111.145 0 111.845 559.045 ;
 RECT 112.945 0 113.645 559.045 ;
 RECT 114.745 0 115.445 559.045 ;
 RECT 116.545 0 117.245 559.045 ;
 RECT 118.345 0 119.045 559.045 ;
 RECT 120.145 0 120.845 559.045 ;
 RECT 121.945 0 122.645 559.045 ;
 RECT 123.745 0 124.445 559.045 ;
 RECT 125.545 0 126.295 559.045 ;
 RECT 127.395 0 129.05 559.045 ;
 RECT 130.15 0 133.885 559.045 ;
 RECT 137.275 0 137.605 559.045 ;
 RECT 139.935 0 140.265 559.045 ;
 RECT 142.595 0 142.925 559.045 ;
 RECT 145.255 0 145.585 559.045 ;
 RECT 147.915 0 148.245 559.045 ;
 RECT 150.575 0 150.905 559.045 ;
 RECT 153.235 0 153.565 559.045 ;
 RECT 155.895 0 156.225 559.045 ;
 RECT 159.615 0 159.945 559.045 ;
 RECT 162.275 0 162.605 559.045 ;
 RECT 164.935 0 165.265 559.045 ;
 RECT 167.595 0 167.925 559.045 ;
 RECT 170.255 0 170.585 559.045 ;
 RECT 172.915 0 173.245 559.045 ;
 RECT 175.575 0 175.905 559.045 ;
 RECT 178.235 0 178.565 559.045 ;
 RECT 181.955 0 182.34 559.045 ;
 END
END S013LLLPSP_X256Y8D8
END LIBRARY
