//**********************************************************************************************
// 16-bit carry look-ahead adder
// Version 0.1
// Modified 17.02.2004
// Designed by Ruslan Lepetenok
// Modified 26.05.12 (Verilog version)
//**********************************************************************************************

`timescale 1 ns / 1 ns

module CLA16B(a_in, b_in, c_in, s_out, c_out);
   input [15:0]  a_in;
   input [15:0]  b_in;
   input         c_in;
   output [15:0] s_out;
   output        c_out;
   
   logic [15:0]   G;
   logic [15:0]   P;
   logic [15:0]   Co;
   
   assign G = a_in & b_in;
   assign P = a_in | b_in;
   
   // Carry generation
   assign Co[0] = G[0] | (P[0] & c_in);
   
   assign Co[1] = G[1] | (P[1] & G[0]) | (P[1] & P[0] & c_in);
   
   assign Co[2] = G[2] | (P[2] & G[1]) | (P[2] & P[1] & G[0]) | (P[2] & P[1] & P[0] & c_in);
   
   assign Co[3] = G[3] | (P[3] & G[2]) | (P[3] & P[2] & G[1]) | (P[3] & P[2] & P[1] & G[0]) | (P[3] & P[2] & P[1] & P[0] & c_in);
   //
   
   assign Co[4] = G[4] | (P[4] & G[3]) | (P[4] & P[3] & G[2]) | (P[4] & P[3] & P[2] & G[1]) | (P[4] & P[3] & P[2] & P[1] & G[0]) | (P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[5] = G[5] | (P[5] & G[4]) | (P[5] & P[4] & G[3]) | (P[5] & P[4] & P[3] & G[2]) | (P[5] & P[4] & P[3] & P[2] & G[1]) | (P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[6] = G[6] | (P[6] & G[5]) | (P[6] & P[5] & G[4]) | (P[6] & P[5] & P[4] & G[3]) | (P[6] & P[5] & P[4] & P[3] & G[2]) | (P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[7] = G[7] | (P[7] & G[6]) | (P[7] & P[6] & G[5]) | (P[7] & P[6] & P[5] & G[4]) | (P[7] & P[6] & P[5] & P[4] & G[3]) | (P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   //		 
   assign Co[8] = G[8] | (P[8] & G[7]) | (P[8] & P[7] & G[6]) | (P[8] & P[7] & P[6] & G[5]) | (P[8] & P[7] & P[6] & P[5] & G[4]) | (P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[9] = G[9] | (P[9] & G[8]) | (P[9] & P[8] & G[7]) | (P[9] & P[8] & P[7] & G[6]) | (P[9] & P[8] & P[7] & P[6] & G[5]) | (P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[10] = G[10] | (P[10] & G[9]) | (P[10] & P[9] & G[8]) | (P[10] & P[9] & P[8] & G[7]) | (P[10] & P[9] & P[8] & P[7] & G[6]) | (P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[11] = G[11] | (P[11] & G[10]) | (P[11] & P[10] & G[9]) | (P[11] & P[10] & P[9] & G[8]) | (P[11] & P[10] & P[9] & P[8] & G[7]) | (P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[12] = G[12] | (P[12] & G[11]) | (P[12] & P[11] & G[10]) | (P[12] & P[11] & P[10] & G[9]) | (P[12] & P[11] & P[10] & P[9] & G[8]) | (P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[13] = G[13] | (P[13] & G[12]) | (P[13] & P[12] & G[11]) | (P[13] & P[12] & P[11] & G[10]) | (P[13] & P[12] & P[11] & P[10] & G[9]) | (P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[14] = G[14] | (P[14] & G[13]) | (P[14] & P[13] & G[12]) | (P[14] & P[13] & P[12] & G[11]) | (P[14] & P[13] & P[12] & P[11] & G[10]) | (P[14] & P[13] & P[12] & P[11] & P[10] & G[9]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   assign Co[15] = G[15] | (P[15] & G[14]) | (P[15] & P[14] & G[13]) | (P[15] & P[14] & P[13] & G[12]) | (P[15] & P[14] & P[13] & P[12] & G[11]) | (P[15] & P[14] & P[13] & P[12] & P[11] & G[10]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & G[9]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & G[8]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & G[7]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & G[6]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & G[5]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & G[4]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & G[3]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[15] & P[14] & P[13] & P[12] & P[11] & P[10] & P[9] & P[8] & P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & c_in);
   
   // Sum generation
   assign s_out[0] = a_in[0] ^ b_in[0] ^ c_in;

      
      assign s_out[15:1] = a_in[15:1] ^ b_in[15:1] ^ Co[14:0];
      
      assign c_out = Co[15]; // Conversion problem was fixed
      
endmodule // CLA16B

// For the purpose of test only (generates wrong result)
// c_out <= Co(Co'high-1);
// For the purpose of test only
