

.SUBCKT inv A VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS N15LL W=nw L=nl m=1
MM1 Y A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS


.SUBCKT STRAP_CELL WL VSS
MN0 VSS WL VSS VSS N15LL W=0.075u L=0.175u m=1
MN1 VSS WL VSS VSS N15LL W=0.075u L=0.175u m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_YMUXB BL BLX DBA DBAX DIN DINX VDDP VSS YS
*.PININFO DIN:I DINX:I YS:I BL:B BLX:B DBA:B DBAX:B VDD:B VSS:B
XI7 YS VDDP VSS net81 / inv pl=130n pw=800n nl=130n nw=800n
XI4 net81 VDDP VSS SL / inv pl=130.00n pw=1.2u nl=130.00n nw=800.0n
MN0 BL DINX net58 VSS N15LL W=2.8u L=130.00n m=1
MN2 BLX DIN net58 VSS N15LL W=2.8u L=130.00n m=1
MN3 net58 SL VSS VSS N15LL W=2.8u L=130.00n m=1
MP0 BL SL VDDP VDDP P15LL W=1u L=130.00n m=1
MP1 BLX SL VDDP VDDP P15LL W=1u L=130.00n m=1
MP2 BL SL BLX VDDP P15LL W=1u L=130.00n m=1
MP3 DBA net81 BL VDDP P15LL W=1.2u L=130.00n m=1
MP4 DBAX net81 BLX VDDP P15LL W=1.2u L=130.00n m=1
.ENDS


.SUBCKT nor2 A B VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 Y B VSS VSS N15LL W=nw L=nl m=1
MM2 Y A VSS VSS N15LL W=nw L=nl m=1
MM1 Y B net35 VDDP P15LL W=pw L=pl m=1
MM0 net35 A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS


.SUBCKT S013EELPSP_delayline_2p4 VDDP VSS Vin Vout
*.PININFO Vin:I Vout:O VDD:B VSS:B
XI275 Vin VDDP VSS net145 / inv pl=130.00n pw=2u nl=130.00n nw=1u
MM0 Vout net145 VDDP VDDP P15LL W=4u L=130.00n m=1
MM1 Vout net145 VSS VSS N15LL W=2u L=130.00n m=1
.ENDS



.SUBCKT buffer_split_right0_mode A SM VDDP VSS Y
*.PININFO A:I SM:I Y:O VDD:B VSS:B
XI143 A net0861 SM VDDP VSS Y / MUX2
XI142 VDDP VSS A net0861 / S013EELPSP_delayline_2p4
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_Logic_OPDEC OP[1] OP[0] S[3] S[2] S[1] S[0] VDDP VSS
*.PININFO OP[1]:I OP[0]:I S[3]:O S[2]:O S[1]:O S[0]:O VDD:B VSS:B
XI34 A BX VDDP VSS S[2] / nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI35 A B VDDP VSS S[0] / nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI27 AX BX VDDP VSS S[3] / nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI31 AX B VDDP VSS S[1] / nand2 pl=130.0n pw=800.0n nl=130.0n nw=800.0n
XI33 BX VDDP VSS B / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI32 AX VDDP VSS A / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI1 OP[1] VDDP VSS BX / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI0 OP[0] VDDP VSS AX / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_FIXDL EMCLK IN OP[1] OP[0] VDDP VSS prc
*.PININFO IN:I OP[1]:I OP[0]:I EMCLK:O prc:O VDD:B VSS:B
XI22 VDDP VSS net36 net37 / S013EELPSP_LEAFCELL_delay100p
XI20 VDDP VSS net40 net36 / S013EELPSP_LEAFCELL_delay100p
XI19 VDDP VSS net44 net40 / S013EELPSP_LEAFCELL_delay100p
XI25 net37 SX[3] S[3] VDDP VSS EMCLK / tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI126 net40 SX[1] S[1] VDDP VSS EMCLK / tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI24 net36 SX[2] S[2] VDDP VSS EMCLK / tgate pl=130.00n pw=5u nl=130.00n nw=5u
XI144 net44 SX[0] S[0] VDDP VSS EMCLK / tgate pl=130.00n pw=4u nl=130.00n nw=4u
XI136 IN VDDP VSS prc / inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
XI137 prc VDDP VSS net44 / inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
XI3[3] S[3] VDDP VSS SX[3] / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[2] S[2] VDDP VSS SX[2] / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[1] S[1] VDDP VSS SX[1] / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI3[0] S[0] VDDP VSS SX[0] / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI0 OP[1] OP[0] S[3] S[2] S[1] S[0] VDDP VSS / S013EELPSP_LEAFCELL_Logic_OPDEC
.ENDS



.SUBCKT S013EELPSP_LEAFCELL_CLKDRV_mode_V1 ACTRCLK ACTRCLKX ACTRCLKX_right  ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right DCTRCLK_right EMCLK  FB_right INTCLKX INTCLKX_right S[1] S[0] SACK1 SACK1_right SACK4 SACK4_right  SM VDDP VMINE VSS WE WEN WE_right
*.PININFO CEN:I CLK:I FB_right:I S[1]:I S[0]:I SM:I VMINE:I WEN:I ACTRCLK:O 
*.PININFO ACTRCLKX:O ACTRCLKX_right:O ACTRCLK_right:O DCTRCLK:O DCTRCLKX:O 
*.PININFO DCTRCLKX_right:O DCTRCLK_right:O EMCLK:O INTCLKX:O INTCLKX_right:O 
*.PININFO SACK1:O SACK1_right:O SACK4:O SACK4_right:O WE:O WE_right:O VDD:B 
*.PININFO VSS:B
XI215 WE SM VDDP VSS WE_right / buffer_split_right0_mode
XI197 CLKLATCH SM VDDP VSS net0257 / buffer_split_right0_mode
XI173 EMCLK CLKLATCH S[1] S[0] VDDP VSS prc_right / S013EELPSP_LEAFCELL_FIXDL
XI134 TESTB net285 VDDP VSS net168 / nand2 pl=130n pw=3u nl=130n nw=3u
XI175 net0397 net0411 VDDP VSS net0194 / nor2 pl=130n pw=6u nl=130n nw=3u
XI174 net0342 net0397 VDDP VSS net0199 / nor2 pl=130n pw=5u nl=130n nw=5u
XI128 CENINT CLK_BUF VDDP VSS net173 / nor2 pl=130n pw=2u nl=130n nw=1.0u
XI143 net337 PRESACK1 VDDP VSS net178 / nor2 pl=130n pw=5u nl=130n nw=5u
XI151 PRESACK1 CLKD VDDP VSS net183 / nor2 pl=130n pw=6u nl=130n nw=3u
MM2 net186 CEN net190 VSS N15LL W=2u L=130.00n m=1
MM3 net190 net261 VSS VSS N15LL W=2u L=130.00n m=1
MM5 CLKLATCH CLK_BUF net198 VSS N15LL W=20u L=130.00n m=1
MM6 net198 net0214 VSS VSS N15LL W=20u L=130.00n m=1
MM1 net186 CEN net205 VDDP P15LL W=2u L=130.00n m=1
MM0 net205 CLK_BUF VDDP VDDP P15LL W=2u L=130.00n m=1
MM11 CLKLATCH CLK_BUF up2 VDDP P15LL W=8.0u L=130.00n m=1
MM4 CLKLATCH net168 VDDP VDDP P15LL W=10u L=130.00n m=1
MM7 FB_right prc_right VDDP VDDP P15LL W=4.8u L=130.00n m=1
MM10 up2 TESTB VDDP VDDP P15LL W=8.0u L=130.00n m=1
XI114 net241 ACTRCLKX ACTRCLK VDDP VSS WENLATCH / tgate pl=130n pw=2u nl=130n  nw=2u
XI212 net0397 VDDP VSS net0344 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI214 net0352 VDDP VSS net0227 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI209 CLK VDDP VSS net0222 / inv pl=130n pw=2.0000u nl=130n nw=1.2u
XI210 net0222 VDDP VSS CLK_BUF / inv pl=130n pw=4u nl=130n nw=2.4u
XI169 VMINE VDDP VSS TESTB / inv pl=130n pw=2.0u nl=130n nw=1.0u
XI188 net0397 VDDP VSS INTCLKX_right / inv pl=130n pw=10u nl=130n nw=10u
XI186 net0194 VDDP VSS SACK4_right / inv pl=130n pw=10u nl=130n nw=5u
XI177 net0257 VDDP VSS net0397 / inv pl=130.00n pw=20u nl=130.00n nw=10u
XI183 net0199 VDDP VSS DCTRCLK_right / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI182 net0199 VDDP VSS net0326 / inv pl=130.00n pw=6u nl=130.00n nw=6u
XI184 net0348 VDDP VSS net0330 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI179 net0199 VDDP VSS ACTRCLK_right / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI178 net0397 VDDP VSS net0257 / inv pl=200.0n pw=250.00n nl=1u nw=250.00n
XI189 net0350 VDDP VSS net0342 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI185 net0330 VDDP VSS net0411 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI176 net0397 VDDP VSS net0350 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI181 net0326 VDDP VSS DCTRCLKX_right / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI180 ACTRCLK_right VDDP VSS ACTRCLKX_right / inv pl=130.00n pw=10u nl=130.00n  nw=5u
XI110 WEN VDDP VSS net237 / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI211 net0344 VDDP VSS net0348 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI112 net237 VDDP VSS net241 / inv pl=300n pw=2u nl=300n nw=2u
XI115 WENLATCH VDDP VSS net245 / inv pl=130n pw=2u nl=130n nw=2u
XI116 net245 VDDP VSS WENLATCH / inv pl=300n pw=250.00n nl=600n nw=250.00n
XI208 net281 VDDP VSS net0214 / inv pl=130n pw=6u nl=130n nw=3u
XI117 net245 VDDP VSS net253 / inv pl=130n pw=6u nl=130n nw=4u
XI118 net253 VDDP VSS WE / inv pl=130n pw=10u nl=130n nw=5u
XI125 CLK_BUF VDDP VSS net261 / inv pl=130n pw=800.0n nl=130n nw=800.0n
XI126 net186 VDDP VSS CENINT / inv pl=130n pw=1.6u nl=130n nw=800.0n
XI127 CENINT VDDP VSS net186 / inv pl=300n pw=250.00n nl=600n nw=250.00n
XI166 PRESACK1 VDDP VSS net273 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI129 net173 VDDP VSS net277 / inv pl=130n pw=2u nl=130n nw=1.0u
XI130 net0334 VDDP VSS net281 / inv pl=130n pw=4u nl=130n nw=2u
XI207 net277 VDDP VSS net0334 / inv pl=130n pw=4u nl=130n nw=2u
XI133 FB_right VDDP VSS net285 / inv pl=130n pw=1.6u nl=130n nw=1.6u
XI141 CLKLATCH VDDP VSS PRESACK1 / inv pl=130.00n pw=20u nl=130.00n nw=10u
XI142 PRESACK1 VDDP VSS CLKLATCH / inv pl=200.0n pw=250.00n nl=1u nw=250.00n
XI187 net0397 VDDP VSS SACK1_right / inv pl=130n pw=10u nl=130n nw=5u
XI144 net178 VDDP VSS ACTRCLK / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI145 ACTRCLK VDDP VSS ACTRCLKX / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI146 net309 VDDP VSS DCTRCLKX / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI147 net178 VDDP VSS net309 / inv pl=130.00n pw=6u nl=130.00n nw=6u
XI148 net178 VDDP VSS DCTRCLK / inv pl=130.00n pw=10u nl=130.00n nw=5u
XI149 net0227 VDDP VSS net317 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI150 net317 VDDP VSS CLKD / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI152 net183 VDDP VSS SACK4 / inv pl=130n pw=10u nl=130n nw=5u
XI153 PRESACK1 VDDP VSS SACK1 / inv pl=130n pw=10u nl=130n nw=5u
XI156 PRESACK1 VDDP VSS INTCLKX / inv pl=130n pw=10u nl=130n nw=10u
XI213 PRESACK1 VDDP VSS net0352 / inv pl=400n pw=800.0n nl=400n nw=800.0n
XI167 net273 VDDP VSS net337 / inv pl=400n pw=800.0n nl=400n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_ESDA13 A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2]  A[1] A[0] CEN CLK S[1] S[0] VDDP VSS WEN
*.PININFO A[10]:I A[9]:I A[8]:I A[7]:I A[6]:I A[5]:I A[4]:I A[3]:I A[2]:I 
*.PININFO A[1]:I A[0]:I CEN:I CLK:I S[1]:I S[0]:I WEN:I VDD:B VSS:B
MM0 A[10] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN29 A[5] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN30 A[6] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN31 A[8] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN32 A[7] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM1 A[9] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN28 WEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 S[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM13 S[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN7 A[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN6 A[2] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN5 A[4] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN4 A[3] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 CEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN2 A[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN0 CLK VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP29 A[5] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP30 A[6] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP31 A[8] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP32 A[7] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP28 WEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM2 A[10] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM3 A[9] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 S[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM15 S[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP7 A[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP6 A[2] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP5 A[4] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP4 A[3] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 CEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP2 A[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP0 CLK VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_ESDA14 A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2]  A[1] A[0] CEN CLK S[1] S[0] VDDP VSS WEN
*.PININFO A[10]:I A[9]:I A[8]:I A[7]:I A[6]:I A[5]:I A[4]:I A[3]:I A[2]:I 
*.PININFO A[1]:I A[0]:I CEN:I CLK:I S[1]:I S[0]:I WEN:I VDD:B VSS:B
MM0 A[10] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM1110 A[11] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN29 A[5] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN30 A[6] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN31 A[8] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN32 A[7] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM1 A[9] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN28 WEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 S[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM13 S[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN7 A[1] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN6 A[2] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN5 A[4] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN4 A[3] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 CEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN2 A[0] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN0 CLK VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP29 A[5] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP30 A[6] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP31 A[8] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP32 A[7] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP28 WEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM2 A[10] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1112 A[11] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM3 A[9] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 S[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM15 S[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP7 A[1] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP6 A[2] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP5 A[4] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP4 A[3] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 CEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP2 A[0] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP0 CLK VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_PXA A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] RDE  VDDP VSS
*.PININFO A[0]:I A[1]:I CLK:I CLKX:I RDE:I PX[3]:O PX[2]:O PX[1]:O PX[0]:O 
*.PININFO VDD:B VSS:B
XI19 net83 CLKX CLK VDDP VSS net59 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI18 net88 CLKX CLK VDDP VSS net65 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI14 net93 CLKX CLK VDDP VSS net71 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI10 net98 CLKX CLK VDDP VSS ALATCH / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI21 AinX[0] Ain[1] VDDP VSS net83 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI20 Ain[0] Ain[1] VDDP VSS net88 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI15 Ain[0] AinX[1] VDDP VSS net93 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI9 AinX[0] AinX[1] VDDP VSS net98 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI62 A[0] VDDP VSS net100 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI25 net59 VDDP VSS PX[2] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI24 PX[2] VDDP VSS net59 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 PX[3] VDDP VSS net65 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI22 net65 VDDP VSS PX[3] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI17 net71 VDDP VSS PX[1] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI16 PX[1] VDDP VSS net71 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI12 PX[0] VDDP VSS ALATCH / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI11 ALATCH VDDP VSS PX[0] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI3 AinX[1] VDDP VSS Ain[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI2 A[1] VDDP VSS AinX[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI1 net100 RDE VDDP VSS Ain[0] / nor2 pl=130.00n pw=2u nl=130.00n nw=1u
XI0 A[0] RDE VDDP VSS AinX[0] / nor2 pl=130.00n pw=1.5u nl=130.00n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_PX4 A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDDP  VSS
*.PININFO A[0]:I A[1]:I CLK:I CLKX:I PX[3]:O PX[2]:O PX[1]:O PX[0]:O VDD:B 
*.PININFO VSS:B
XI19 net94 CLKX CLK VDDP VSS net70 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI18 net99 CLKX CLK VDDP VSS net76 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI14 net104 CLKX CLK VDDP VSS net82 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI10 net109 CLKX CLK VDDP VSS net88 / tgate pl=130.00n pw=3u nl=130.00n nw=3u
XI21 AinX[0] Ain[1] VDDP VSS net94 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI20 Ain[0] Ain[1] VDDP VSS net99 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI15 Ain[0] AinX[1] VDDP VSS net104 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI9 AinX[0] AinX[1] VDDP VSS net109 / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI25 net70 VDDP VSS PX[2] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI24 PX[2] VDDP VSS net70 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 PX[3] VDDP VSS net76 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI22 net76 VDDP VSS PX[3] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI17 net82 VDDP VSS PX[1] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI16 PX[1] VDDP VSS net82 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI12 PX[0] VDDP VSS net88 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI11 net88 VDDP VSS PX[0] / inv pl=130.00n pw=7u nl=130.00n nw=2u
XI3 AinX[1] VDDP VSS Ain[1] / inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI2 A[1] VDDP VSS AinX[1] / inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI1 AinX[0] VDDP VSS Ain[0] / inv pl=130.00n pw=2u nl=130.00n nw=1.4u
XI0 A[0] VDDP VSS AinX[0] / inv pl=130.00n pw=2u nl=130.00n nw=1.4u
.ENDS

.SUBCKT nand3 A B C VDDP VSS Y pw=1u pl=180.0n nw=1u nl=180.0n
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM6 net29 C VSS VSS N15LL W=nw L=nl m=1
MM5 net33 B net29 VSS N15LL W=nw L=nl m=1
MM4 Y A net33 VSS N15LL W=nw L=nl m=1
MM3 Y A VDDP VDDP P15LL W=pw L=pl m=1
MM2 Y B VDDP VDDP P15LL W=pw L=pl m=1
MM1 Y C VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_FPREDEC_YX A[0] A[1] CLK CLKX FCKX[3] FCKX[2]  FCKX[1] FCKX[0] VDDP VSS WLCKX
*.PININFO A[0]:I A[1]:I CLK:I CLKX:I WLCKX:I FCKX[3]:O FCKX[2]:O FCKX[1]:O 
*.PININFO FCKX[0]:O VDD:B VSS:B
XI187 Ain[0] AinX[1] VDDP VSS net221 / nand2 pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI196 AinX[0] Ain[1] VDDP VSS net227 / nand2 pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI195 Ain[0] Ain[1] VDDP VSS net233 / nand2 pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI133 AinX[0] AinX[1] VDDP VSS net268 / nand2 pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI191 net270 WLCKX VDDP VSS net135 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI192 net326 WLCKX VDDP VSS net140 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI185 net274 WLCKX VDDP VSS net145 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI183 net314 WLCKX VDDP VSS net170 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI186 net221 CLKX CLK VDDP VSS net175 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI194 net227 CLKX CLK VDDP VSS net181 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI193 net233 CLKX CLK VDDP VSS net187 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI134 net268 CLKX CLK VDDP VSS FALATCH / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI229 net366 VDDP VSS net270 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI228 net390 VDDP VSS net274 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI188 net145 VDDP VSS FCKX[1] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI189 net390 VDDP VSS net175 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI235 A[0] VDDP VSS net302 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI199 net135 VDDP VSS FCKX[3] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI201 net410 VDDP VSS net181 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI227 net359 VDDP VSS net314 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI230 net410 VDDP VSS net326 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI136 net359 VDDP VSS FALATCH / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI135 FALATCH VDDP VSS net359 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI197 net187 VDDP VSS net366 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI184 net170 VDDP VSS FCKX[0] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI190 net175 VDDP VSS net390 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI198 net366 VDDP VSS net187 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI200 net140 VDDP VSS FCKX[2] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI202 net181 VDDP VSS net410 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI236 A[1] VDDP VSS net414 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI137 Ain[1] VDDP VSS AinX[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI2 net414 VDDP VSS Ain[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI132 Ain[0] VDDP VSS AinX[0] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI0 net302 VDDP VSS Ain[0] / inv pl=130.00n pw=2u nl=130.00n nw=1u
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_FPREDEC A[0] A[1] A[2] CLK CLKX FCKX[7] FCKX[6]  FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] VDDP VSS WLCKX
*.PININFO A[0]:I A[1]:I A[2]:I CLK:I CLKX:I WLCKX:I FCKX[7]:O FCKX[6]:O 
*.PININFO FCKX[5]:O FCKX[4]:O FCKX[3]:O FCKX[2]:O FCKX[1]:O FCKX[0]:O VDD:B 
*.PININFO VSS:B
XI191 net270 WLCKX VDDP VSS net135 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI192 net326 WLCKX VDDP VSS net140 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI185 net274 WLCKX VDDP VSS net145 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI203 net286 WLCKX VDDP VSS net150 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI204 net282 WLCKX VDDP VSS net155 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI205 net318 WLCKX VDDP VSS net160 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI206 net278 WLCKX VDDP VSS net165 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI183 net314 WLCKX VDDP VSS net170 / nor2 pl=130.0n pw=4u nl=130.0n nw=2u
XI186 net221 CLKX CLK VDDP VSS net175 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI194 net227 CLKX CLK VDDP VSS net181 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI193 net233 CLKX CLK VDDP VSS net187 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI207 net239 CLKX CLK VDDP VSS net193 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI208 net245 CLKX CLK VDDP VSS net199 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI209 net257 CLKX CLK VDDP VSS net205 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI210 net251 CLKX CLK VDDP VSS net211 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI134 net268 CLKX CLK VDDP VSS net0730 / tgate pl=130.00n pw=1.5u nl=130.00n  nw=1.5u
XI187 Ain[0] AinX[1] AinX[2] VDDP VSS net221 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI196 AinX[0] Ain[1] AinX[2] VDDP VSS net227 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI195 Ain[0] Ain[1] AinX[2] VDDP VSS net233 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI211 AinX[0] Ain[1] Ain[2] VDDP VSS net239 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI212 Ain[0] Ain[1] Ain[2] VDDP VSS net245 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI214 AinX[0] AinX[1] Ain[2] VDDP VSS net251 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI213 Ain[0] AinX[1] Ain[2] VDDP VSS net257 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI133 AinX[0] AinX[1] AinX[2] VDDP VSS net268 / nand3 pl=130.00n pw=1.5u  nl=130.00n nw=1.5u
XI229 net0346 VDDP VSS net270 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI228 net0334 VDDP VSS net274 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI234 net0182 VDDP VSS net278 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI232 net0370 VDDP VSS net282 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI231 net0277 VDDP VSS net286 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI188 net145 VDDP VSS FCKX[1] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI189 net0334 VDDP VSS net175 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI237 A[2] VDDP VSS net298 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI235 A[0] VDDP VSS net302 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI199 net135 VDDP VSS FCKX[3] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI201 net0318 VDDP VSS net181 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI227 net359 VDDP VSS net314 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI233 net0342 VDDP VSS net318 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI220 net199 VDDP VSS net0370 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI230 net0318 VDDP VSS net326 / inv pl=130.00n pw=2.2u nl=130.00n nw=2.2u
XI82 net298 VDDP VSS Ain[2] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI215 net193 VDDP VSS net0277 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI217 net150 VDDP VSS FCKX[6] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI216 net0277 VDDP VSS net193 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI218 net155 VDDP VSS FCKX[7] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI138 Ain[2] VDDP VSS AinX[2] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI136 net359 VDDP VSS net0730 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI135 net0730 VDDP VSS net359 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI219 net0370 VDDP VSS net199 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI197 net187 VDDP VSS net0346 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI221 net205 VDDP VSS net0342 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI223 net160 VDDP VSS FCKX[5] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI224 net165 VDDP VSS FCKX[4] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI184 net170 VDDP VSS FCKX[0] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI225 net0182 VDDP VSS net211 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI190 net175 VDDP VSS net0334 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI222 net0342 VDDP VSS net205 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI226 net211 VDDP VSS net0182 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI198 net0346 VDDP VSS net187 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI200 net140 VDDP VSS FCKX[2] / inv pl=130.00n pw=5u nl=130.00n nw=5u
XI202 net181 VDDP VSS net0318 / inv pl=130.00n pw=1.1u nl=130.00n nw=1.1u
XI236 A[1] VDDP VSS net414 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI137 Ain[1] VDDP VSS AinX[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI2 net414 VDDP VSS Ain[1] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI132 Ain[0] VDDP VSS AinX[0] / inv pl=130.00n pw=2u nl=130.00n nw=1u
XI0 net302 VDDP VSS Ain[0] / inv pl=130.00n pw=2u nl=130.00n nw=1u
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_TieL_S TieL VDDP VSS
*.PININFO TieL:O VDD:B VSS:B
MN18 TieL net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 net15 net15 VDDP VDDP P15LL W=1.6u L=130.00n m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_TieH_S Tie_high VDDP VSS
*.PININFO Tie_high:O VDD:B VSS:B
MN18 net15 net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 Tie_high net15 VDDP VDDP P15LL W=3u L=130.00n m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_STWL_DEC EMCLK STWL VDDP VSS
*.PININFO EMCLK:I STWL:O VDD:B VSS:B
MP9 A T_HIGH VDDP VDDP P15LL W=800.0n L=130.00n m=1
MP18 net61 net61 VDDP VDDP P15LL W=800.0n L=130.00n m=1
MM4 T_HIGH net77 VDDP VDDP P15LL W=2u L=130.00n m=1
MM0 STWL C VDDP VDDP P15LL W=5u L=130.00n m=1
MM5 net77 net77 VSS VSS N15LL W=800.0n L=130.00n m=1
MN18 T_LOW net61 VSS VSS N15LL W=1u L=130.00n m=1
MM1 STWL C VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS C / inv pl=130.00n pw=3u nl=130.00n nw=3u
XI8 A VDDP VSS B / inv pl=130.00n pw=1u nl=130.00n nw=1u
XI114 A T_HIGH T_LOW VDDP VSS EMCLK / tgate pl=130.00n pw=800.0n nl=130.00n  nw=1.2u
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_DischargeCells DUM_BL EMCLK S[2] S[1] S[0] VDDP VSS
*.PININFO EMCLK:I S[2]:I S[1]:I S[0]:I DUM_BL:B VDD:B VSS:B
MN6 net30 S[2] VSS VSS NPD W=220.000n L=130.000n m=8
MN5 net34 S[1] VSS VSS NPD W=220.000n L=130.000n m=4
MN2 net38 S[0] VSS VSS NPD W=220.000n L=130.000n m=4
MN1 net42 VDDP VSS VSS NPD W=220.000n L=130.000n m=4
MN16 DUM_BL EMCLK net42 VSS NPG W=150.000n L=175.00n m=4
MN7 DUM_BL EMCLK net30 VSS NPG W=150.000n L=175.00n m=8
MN4 DUM_BL EMCLK net34 VSS NPG W=150.000n L=175.00n m=4
MN3 DUM_BL EMCLK net38 VSS NPG W=150.000n L=175.00n m=4
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_OPDEC OP[1] OP[0] S[2] S[1] S[0] VDDP VSS
*.PININFO OP[1]:I OP[0]:I S[2]:O S[1]:O S[0]:O VDD:B VSS:B
XI12 AX BX VDDP VSS S[2] / nor2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI6 AX BX VDDP VSS S[0] / nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI7 BX VDDP VSS S[1] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI1 OP[1] VDDP VSS BX / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI0 OP[0] VDDP VSS AX / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_SOP DBL_right EMCLK S[2] S[3] STWL_right VDDP VSS
*.PININFO EMCLK:I S[2]:I S[3]:I DBL_right:O STWL_right:O VDD:B VSS:B
XI16 TieLS VDDP VSS / S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013EELPSP_LEAFCELL_TieH_S
MM0 S[2] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 S[3] VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 S[2] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 S[3] VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013EELPSP_LEAFCELL_DischargeCells
XI21 S[3] S[2] OP[2] OP[1] OP[0] VDDP VSS / S013EELPSP_LEAFCELL_OPDEC
.ENDS
.SUBCKT S013EELPSP_SOP00 DBL_right EMCLK STWL_right VDDP VSS
*.PININFO EMCLK:I S[2]:I S[3]:I DBL_right:O STWL_right:O VDD:B VSS:B
XI16 TieLS VDDP VSS / S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013EELPSP_LEAFCELL_TieH_S
MM0 TieLS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 TieLS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 TieLS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 TieLS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013EELPSP_LEAFCELL_DischargeCells
XI21 TieLS TieLS OP[2] OP[1] OP[0] VDDP VSS / S013EELPSP_LEAFCELL_OPDEC
.ENDS
.SUBCKT S013EELPSP_SOP01 DBL_right EMCLK STWL_right VDDP VSS
*.PININFO EMCLK:I TieHS:I TieLS:I DBL_right:O STWL_right:O VDD:B VSS:B
XI16 TieLS VDDP VSS / S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013EELPSP_LEAFCELL_TieH_S
MM0 TieHS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 TieLS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 TieHS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 TieLS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013EELPSP_LEAFCELL_DischargeCells
XI21 TieLS TieHS OP[2] OP[1] OP[0] VDDP VSS / S013EELPSP_LEAFCELL_OPDEC
.ENDS
SUBCKT S013EELPSP_SOP10 DBL_right EMCLK  STWL_right VDDP VSS
*.PININFO EMCLK:I TieLS:I TieHS:I DBL_right:O STWL_right:O VDD:B VSS:B
XI16 TieLS VDDP VSS / S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013EELPSP_LEAFCELL_TieH_S
MM0 TieLS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 TieHS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 TieLS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 TieHS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013EELPSP_LEAFCELL_DischargeCells
XI21 TieHS TieLS OP[2] OP[1] OP[0] VDDP VSS / S013EELPSP_LEAFCELL_OPDEC
.ENDS
.SUBCKT S013EELPSP_SOP11 DBL_right EMCLK STWL_right VDDP VSS
*.PININFO EMCLK:I TieHS:I TieHS:I DBL_right:O STWL_right:O VDD:B VSS:B
XI16 TieLS VDDP VSS / S013EELPSP_LEAFCELL_TieL_S
XI17 TieHS VDDP VSS / S013EELPSP_LEAFCELL_TieH_S
MM0 TieHS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM11 TieHS VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MM1 TieHS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MM10 TieHS VSS VSS VSS N15LL W=300.0n L=130.00n m=1
XI19 EMCLK STWL_right VDDP VSS / S013EELPSP_LEAFCELL_STWL_DEC
XI18 DBL_right STWL_right OP[2] OP[1] OP[0] VDDP VSS /  S013EELPSP_LEAFCELL_DischargeCells
XI21 TieHS TieHS OP[2] OP[1] OP[0] VDDP VSS / S013EELPSP_LEAFCELL_OPDEC
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_TieH Tie_high VDDP VSS
*.PININFO Tie_high:O VDD:B VSS:B
MN18 net15 net15 VSS VSS N15LL W=2u L=130.00n m=1
MP18 Tie_high net15 VDDP VDDP P15LL W=4u L=130.00n m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_TieL TieL VDDP VSS
*.PININFO TieL:O VDD:B VSS:B
MN18 TieL net15 VSS VSS N15LL W=4u L=130.00n m=1
MP18 net15 net15 VDDP VDDP P15LL W=2u L=130.00n m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_RWL_DEC_left CLK CLKX RDE RWLL VDDP VSS WLCKX
*.PININFO CLK:I CLKX:I RDE:I WLCKX:I RWLL:O VDD:B VSS:B
MP9 net64 net97 VDDP VDDP P15LL W=4u L=130.00n m=1
XI114 net64 net97 net93 VDDP VSS WLCKX / tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI2 net73 CLKX CLK VDDP VSS net69 / tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI3 net77 VDDP VSS net73 / inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI8 RDE VDDP VSS net77 / inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI129 net64 VDDP VSS RWLL / inv pl=130.00n pw=5u nl=130.00n nw=2u
XI1 net93 VDDP VSS net69 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI0 net69 VDDP VSS net93 / inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI24 net93 VDDP VSS net97 / inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_RWL_DEC_right CLK CLKX RDE RWLR VDDP VSS WLCKX
*.PININFO CLK:I CLKX:I RDE:I WLCKX:I RWLR:O VDD:B VSS:B
MP0 net58 net97 VDDP VDDP P15LL W=4u L=130.00n m=1
XI5 net58 net97 net93 VDDP VSS WLCKX / tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI2 net73 CLKX CLK VDDP VSS net69 / tgate pl=130.00n pw=2u nl=130.00n nw=2u
XI3 net77 VDDP VSS net73 / inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI8 RDE VDDP VSS net77 / inv pl=130.00n pw=1u nl=130.00n nw=800.0n
XI7 net58 VDDP VSS RWLR / inv pl=130.00n pw=5u nl=130.00n nw=2u
XI1 net93 VDDP VSS net69 / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI0 net69 VDDP VSS net93 / inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI24 net93 VDDP VSS net97 / inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_FDEC_right FCKX PABC PABCX VDDP VSS WLR
*.PININFO FCKX:I PABC:I PABCX:I WLR:O VDD:B VSS:B
MM2 WLR net46 VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS net46 / inv pl=130.00n pw=3u nl=130.00n nw=3u
XI8 A VDDP VSS B / inv pl=130.00n pw=1u nl=130.00n nw=1u
MM3 WLR net46 VDDP VDDP P15LL W=5u L=130.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
XI114 A PABC PABCX VDDP VSS FCKX / tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_delay100p VDDP VSS in out
*.PININFO in:I out:O VDD:B VSS:B
MM0 net17 in VSS VSS N15LL W=800.0n L=300.00n m=1
MM1 net17 in VDDP VDDP P15LL W=800.0n L=130.00n m=1
XI0 net17 VDDP VSS out / inv pl=130.00n pw=2.8u nl=130.00n nw=1.4u
.ENDS



.SUBCKT MUX2 I0 I1 S VDDP VSS Z
*.PININFO I0:I I1:I S:I Z:O VDD:B VSS:B
XI2 net40 net44 VDDP VSS net030 / nor2 pl=130n pw=2u nl=130n nw=1u
XI8 net030 VDDP VSS Z / inv pl=130n pw=4u nl=130n nw=2u
XI6 net49 VDDP VSS net40 / inv pl=130n pw=2u nl=130n nw=1u
XI4 net54 VDDP VSS net44 / inv pl=130n pw=2u nl=130n nw=1u
XI5 S VDDP VSS net36 / inv pl=130n pw=2u nl=130n nw=1u
XI3 I0 net36 VDDP VSS net54 / nand2 pl=130.0n pw=2u nl=130.0n nw=1u
XI7 I1 S VDDP VSS net49 / nand2 pl=130.0n pw=2u nl=130.0n nw=1u
.ENDS



.SUBCKT nand2 A B VDDP VSS Y pw=1u pl=180.0n nw=1u nl=180.0n
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 Y A net26 VSS N15LL W=nw L=nl m=1
MM0 net26 B VSS VSS N15LL W=nw L=nl m=1
MM2 Y B VDDP VDDP P15LL W=pw L=pl m=1
MM1 Y A VDDP VDDP P15LL W=pw L=pl m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_SA8 DB DBX DOUT VDDP VSS ck1 ck4
*.PININFO ck1:I ck4:I DOUT:O DB:B DBX:B VDD:B VSS:B
MN4 net85 ck3 net94 VSS N15LL W=2u L=130.00n m=1
MN0 DX D net85 VSS N15LL W=6u L=200.0n m=1
MN1 D DX net85 VSS N15LL W=6u L=200.0n m=1
MN3 net94 ck6 VSS VSS N15LL W=2u L=130.00n m=1
MP0 DBX ck6 VDDP VDDP P15LL W=1u L=130.00n m=1
MP1 DB ck6 VDDP VDDP P15LL W=1u L=130.00n m=1
MP2 DB ck6 DBX VDDP P15LL W=1u L=130.00n m=1
MP3 D close DB VDDP P15LL W=2.8u L=130.00n m=1
MP4 DX close DBX VDDP P15LL W=2.8u L=130.00n m=1
MP7 DX D VDDP VDDP P15LL W=1.6u L=200.0n m=1
MP8 D DX VDDP VDDP P15LL W=1.6u L=200.0n m=1
XI53 DX DOUTB VDDP VSS DOUTBB / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI54 DOUTBB D VDDP VSS DOUTB / nand2 pl=130.00n pw=1u nl=130.00n nw=1u
XI74 ck1 ck4 VDDP VSS net137 / nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI73 net156 VDDP VSS ck6 / inv pl=130.00n pw=3.2u nl=130.00n nw=1.6u
XI71 net152 VDDP VSS ck3 / inv pl=130.00n pw=2u nl=130.00n nw=1.0u
XI77 DOUTB VDDP VSS DOUT / inv pl=130.00n pw=3u nl=130.00n nw=1.5u
XI70 ck1 VDDP VSS net152 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI72 ck4 VDDP VSS net156 / inv pl=130.00n pw=1.6u nl=130.00n nw=800.0n
XI75 net137 VDDP VSS close / inv pl=130.00n pw=2u nl=130.00n nw=1.0u
.ENDS



.SUBCKT tgate A EN ENX VDDP VSS Y pw=1u pl=180n nw=1u nl=180n
*.PININFO EN:I ENX:I A:B VDD:B VSS:B Y:B
M0 A EN Y VSS N15LL W=nw L=nl m=1
M1 A ENX Y VDDP P15LL W=pw L=pl m=1
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_DATAIN BWEN CLK CLKX D DATA DX VDDP VSS WE
*.PININFO BWEN:I CLK:I CLKX:I DATA:I WE:I D:O DX:O VDD:B VSS:B
XI136 WE net122 VDDP VSS net77 / nand2 pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI4 net142 net126 VDDP VSS net82 / nand2 pl=130.00n pw=800.0n nl=130.00n nw=1u
XI3 net154 net126 VDDP VSS net87 / nand2 pl=130.00n pw=800.0n nl=130.00n nw=1u
XI21 net114 CLKX CLK VDDP VSS BLATCH / tgate pl=130.00n pw=1.4u nl=130.00n  nw=1.4u
XI5 net146 CLKX CLK VDDP VSS DLATCH / tgate pl=130.00n pw=1.4u nl=130.00n  nw=1.4u
XI39 BWEN VDDP VSS net0206 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI37 net0206 VDDP VSS net0207 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI31 net0100 VDDP VSS net0104 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI35 net0207 VDDP VSS net0120 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI34 DATA VDDP VSS net0100 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI30 net0112 VDDP VSS net0108 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI29 net0104 VDDP VSS net0112 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI28 net0108 VDDP VSS net102 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI322 net130 VDDP VSS net106 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI321 net106 VDDP VSS net110 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI320 net110 VDDP VSS net114 / inv pl=130.00n pw=1.4u nl=130.00n nw=1.4u
XI22 net122 VDDP VSS BLATCH / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI23 BLATCH VDDP VSS net122 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI143 net77 VDDP VSS net126 / inv pl=130.00n pw=1.6u nl=130.00n nw=1.0u
XI323 net0146 VDDP VSS net130 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI19 net87 VDDP VSS DX / inv pl=130.00n pw=1.44u nl=130.00n nw=720.00n
XI20 net82 VDDP VSS D / inv pl=130.00n pw=1.44u nl=130.00n nw=720.00n
XI15 net154 VDDP VSS net142 / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI36 net0120 VDDP VSS net0146 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI27 net162 VDDP VSS net146 / inv pl=130.00n pw=1.4u nl=130.00n nw=1.4u
XI9 net154 VDDP VSS DLATCH / inv pl=300.0n pw=250.00n nl=600.0n nw=250.00n
XI7 DLATCH VDDP VSS net154 / inv pl=130.00n pw=1.6u nl=130.00n nw=1.0u
XI25 net102 VDDP VSS net158 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
XI26 net158 VDDP VSS net162 / inv pl=300.0n pw=800.0n nl=300.0n nw=800.0n
.ENDS

.SUBCKT BITCELL B BX VDDC VSS WL1
*.PININFO WL1:I B:B BX:B VDDC:B VSS:B
MM2 BX WL1 BCN VSS NPG W=150.000n L=175.00n m=1
MM3 B WL1 BC VSS NPG W=150.000n L=175.00n m=1
MM0 BCN BC VSS VSS NPD W=220.00n L=130.00n m=1
MM1 BC BCN VSS VSS NPD W=220.00n L=130.00n m=1
MM5 BCN BC VDDC VDDC PL W=160.000n L=150.00n m=1
MM6 BC BCN VDDC VDDC PL W=160.000n L=150.00n m=1
.ENDS


.SUBCKT S013EELPSP_bitcell_STWL B BX VDDC VSS WL
*.PININFO WL:I B:B BX:B VDDC:B VSS:B
MM5 BCN BC VDDC VDDC PL W=160.000n L=150.00n m=1
MM6 BC BCN VDDC VDDC PL W=160.000n L=150.00n m=1
MM0 BCN BC VSS VSS NPD W=220.00n L=130.00n m=1
MM1 BC BCN VSS VSS NPD W=220.00n L=130.00n m=1
MM2 BX WL BCN VSS NPG W=150.000n L=175.00n m=1
MM3 B VSS BC VSS NPG W=150.000n L=175.00n m=1
.ENDS



.SUBCKT S013EELPSP_pcap_st B BX VDDC VSS WL0
*.PININFO WL0:I B:B BX:B VDDC:B VSS:B
MTL1 net42 net51 VDDC VDDC PL W=160.000n L=150.000n m=1
MTL0 net51 net42 VDDC VDDC PL W=160.000n L=150.000n m=1
MTD0 net51 net42 VSS VSS NPD W=220.000n L=130.000n m=1
MTD1 net42 net51 VSS VSS NPD W=220.000n L=130.000n m=1
MTA0 B WL0 net51 VSS NPG W=150.000n L=175.00n m=1
MTA1 BX VSS net42 VSS NPG W=150.000n L=175.00n m=1
.ENDS


.SUBCKT S013EELPSP_pcap B BX VDDC VSS WL
*.PININFO WL:I B:B BX:B VDDC:B VSS:B
MM2 BX WL net034 VSS NPG W=150.000n L=175.00n m=1
MTA1 B WL net27 VSS NPG W=150.000n L=175.00n m=1
MM1 net034 net27 VSS VSS NPD W=220.000n L=130.000n m=1
MTD1 net27 net034 VSS VSS NPD W=220.000n L=130.000n m=1
MM0 net034 net27 VDDC VDDC PL W=160.000n L=150.000n m=1
MTL1 net27 net034 VDDC VDDC PL W=160.000n L=150.000n m=1
.ENDS



.SUBCKT S013EELPSP_pcap_STWL_b STWL[3] STWL[2] STWL[1] STWL[0] VDDC VSS
*.PININFO STWL[3]:I STWL[2]:I STWL[1]:I STWL[0]:I VDDC:B VSS:B
XI4 net029 net027 VDDC VSS STWL[1] / S013EELPSP_pcap
XI6 net14 net019 VDDC VSS STWL[3] / S013EELPSP_pcap
XI5 net14 net019 VDDC VSS STWL[2] / S013EELPSP_pcap
XI3 net029 net027 VDDC VSS STWL[0] / S013EELPSP_pcap
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_XDEC_right FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]  FCKX[2] FCKX[1] FCKX[0] PXA PXB PXC VDDP VSS WLR[7] WLR[6] WLR[5] WLR[4]  WLR[3] WLR[2] WLR[1] WLR[0]
*.PININFO FCKX[7]:I FCKX[6]:I FCKX[5]:I FCKX[4]:I FCKX[3]:I FCKX[2]:I 
*.PININFO FCKX[1]:I FCKX[0]:I PXA:I PXB:I PXC:I WLR[7]:O WLR[6]:O WLR[5]:O 
*.PININFO WLR[4]:O WLR[3]:O WLR[2]:O WLR[1]:O WLR[0]:O VDD:B VSS:B
XI156 PXA PXB PXC VDDP VSS net31 / nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XIFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLR[7] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLR[6] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLR[5] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLR[4] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLR[3] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLR[2] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLR[1] / S013EELPSP_LEAFCELL_FDEC_right
XIFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLR[0] / S013EELPSP_LEAFCELL_FDEC_right
XI111 net31 VDDP VSS PABC / inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_FDEC_left FCKX PABC PABCX VDDP VSS WLL
*.PININFO FCKX:I PABC:I PABCX:I WLL:O VDD:B VSS:B
MM1 WLL C VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS C / inv pl=130.00n pw=3u nl=130.00n nw=3u
XI8 A VDDP VSS B / inv pl=130.00n pw=1u nl=130.00n nw=1u
MM0 WLL C VDDP VDDP P15LL W=5u L=130.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
XI114 A PABC PABCX VDDP VSS FCKX / tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
.ENDS



.SUBCKT S013EELPSP_LEAFCELL_XDEC_left FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]  FCKX[2] FCKX[1] FCKX[0] PXA PXB PXC VDDP VSS WLL[7] WLL[6] WLL[5] WLL[4]  WLL[3] WLL[2] WLL[1] WLL[0]
*.PININFO FCKX[7]:I FCKX[6]:I FCKX[5]:I FCKX[4]:I FCKX[3]:I FCKX[2]:I 
*.PININFO FCKX[1]:I FCKX[0]:I PXA:I PXB:I PXC:I WLL[7]:O WLL[6]:O WLL[5]:O 
*.PININFO WLL[4]:O WLL[3]:O WLL[2]:O WLL[1]:O WLL[0]:O VDD:B VSS:B
XI156 PXA PXB PXC VDDP VSS net31 / nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XIFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLL[7] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLL[6] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLL[5] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLL[4] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLL[3] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLL[2] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLL[1] / S013EELPSP_LEAFCELL_FDEC_left
XIFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLL[0] / S013EELPSP_LEAFCELL_FDEC_left
XI111 net31 VDDP VSS PABC / inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS


/**********YMUX4****************/
.SUBCKT S013EELPSP_LEAFCELL_YMUX4 BL[3] BL[2] BL[1] BL[0] BLX[3] BLX[2] BLX[1]  BLX[0] DB DBX DIN DINX VDDP VSS YS[3] YS[2] YS[1] YS[0]
*.PININFO DIN:I DINX:I YS[3]:I YS[2]:I YS[1]:I YS[0]:I BL[3]:B BL[2]:B BL[1]:B 
*.PININFO BL[0]:B BLX[3]:B BLX[2]:B BLX[1]:B BLX[0]:B DB:B DBX:B VDD:B VSS:B
XI3 BL[3] BLX[3] DB DBX DIN DINX VDDP VSS YS[3] / S013EELPSP_LEAFCELL_YMUXB
XI2 BL[2] BLX[2] DB DBX DIN DINX VDDP VSS YS[2] / S013EELPSP_LEAFCELL_YMUXB
XI1 BL[1] BLX[1] DB DBX DIN DINX VDDP VSS YS[1] / S013EELPSP_LEAFCELL_YMUXB
XI0 BL[0] BLX[0] DB DBX DIN DINX VDDP VSS YS[0] / S013EELPSP_LEAFCELL_YMUXB
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_YMX4SAWR_BW BL[3] BL[2] BL[1] BL[0] BLX[3] BLX[2]  BLX[1] BLX[0] BWEN CLK CLKX DATA DOUT SACK1 SACK4 VDDP VSS WE YX[3] YX[2]  YX[1] YX[0]
*.PININFO BWEN:I CLK:I CLKX:I DATA:I SACK1:I SACK4:I WE:I YX[3]:I YX[2]:I 
*.PININFO YX[1]:I YX[0]:I DOUT:O BL[3]:B BL[2]:B BL[1]:B BL[0]:B BLX[3]:B 
*.PININFO BLX[2]:B BLX[1]:B BLX[0]:B VDD:B VSS:B
XYMUX4 BL[3] BL[2] BL[1] BL[0] BLX[3] BLX[2] BLX[1] BLX[0] DB DBX DIN DINX VDDP  VSS net86[3] net86[2] net86[1] net86[0] / S013EELPSP_LEAFCELL_YMUX4
XSA DB DBX DOUT VDDP VSS SACK1 SACK4 / S013EELPSP_LEAFCELL_SA8
MN1 BWEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 DATA VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP1 BWEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 DATA VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
XI14[3] YX[3] VDDP VSS net86[3] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[2] YX[2] VDDP VSS net86[2] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[1] YX[1] VDDP VSS net86[1] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[0] YX[0] VDDP VSS net86[0] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XIDATAIN BWEN CLK CLKX DIN DATA DINX VDDP VSS WE / S013EELPSP_LEAFCELL_DATAIN
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_Logic_common_mode_Y4 ACTRCLK ACTRCLKX ACTRCLKX_right  ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right DCTRCLK_right EMCLK  FB_right FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0]  FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3]  FCKX_right[2] FCKX_right[1] FCKX_right[0] INTCLKX INTCLKX_right PXA[3]  PXA[2] PXA[1] PXA[0] PXA_right[3] PXA_right[2] PXA_right[1] PXA_right[0]  PXB[3] PXB[2] PXB[1] PXB[0] PXB_right[3] PXB_right[2] PXB_right[1]  PXB_right[0] PXC[3] PXC[2] PXC[1] PXC[0] PXC_right[3] PXC_right[2]  PXC_right[1] PXC_right[0] RDE S[1] S[0] SACK1 SACK1_right SACK4 SACK4_right  SM VDDP VMINE VSS WE WEN WE_right XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2]  XA[1] XA[0] YA[1] YA[0] YX[3] YX[2] YX[1] YX[0] YX_right[3] YX_right[2]  YX_right[1] YX_right[0]
*.PININFO CEN:I CLK:I FB_right:I RDE:I S[1]:I S[0]:I SM:I VMINE:I WEN:I 
*.PININFO XA[8]:I XA[7]:I XA[6]:I XA[5]:I XA[4]:I XA[3]:I XA[2]:I XA[1]:I 
*.PININFO XA[0]:I YA[1]:I YA[0]:I ACTRCLK:O ACTRCLKX:O ACTRCLKX_right:O 
*.PININFO ACTRCLK_right:O DCTRCLK:O DCTRCLKX:O DCTRCLKX_right:O 
*.PININFO DCTRCLK_right:O EMCLK:O FCKX[7]:O FCKX[6]:O FCKX[5]:O FCKX[4]:O 
*.PININFO FCKX[3]:O FCKX[2]:O FCKX[1]:O FCKX[0]:O FCKX_right[7]:O 
*.PININFO FCKX_right[6]:O FCKX_right[5]:O FCKX_right[4]:O FCKX_right[3]:O 
*.PININFO FCKX_right[2]:O FCKX_right[1]:O FCKX_right[0]:O INTCLKX:O 
*.PININFO INTCLKX_right:O PXA[3]:O PXA[2]:O PXA[1]:O PXA[0]:O PXA_right[3]:O 
*.PININFO PXA_right[2]:O PXA_right[1]:O PXA_right[0]:O PXB[3]:O PXB[2]:O 
*.PININFO PXB[1]:O PXB[0]:O PXB_right[3]:O PXB_right[2]:O PXB_right[1]:O 
*.PININFO PXB_right[0]:O PXC[3]:O PXC[2]:O PXC[1]:O PXC[0]:O PXC_right[3]:O 
*.PININFO PXC_right[2]:O PXC_right[1]:O PXC_right[0]:O SACK1:O SACK1_right:O 
*.PININFO SACK4:O SACK4_right:O WE:O WE_right:O YX[3]:O YX[2]:O YX[1]:O 
*.PININFO YX[0]:O YX_right[3]:O YX_right[2]:O YX_right[1]:O YX_right[0]:O 
*.PININFO VDD:B VSS:B
XICLKDRV ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX  DCTRCLKX_right DCTRCLK_right EMCLK FB_right INTCLKX INTCLKX_right S[1] S[0]  SACK1 SACK1_right SACK4 SACK4_right SM VDDP VMINE VSS WE WEN WE_right /  S013EELPSP_LEAFCELL_CLKDRV_mode_V1
XI18 YA[0] YA[1] ACTRCLK_right ACTRCLKX_right YX_right[3] YX_right[2]  YX_right[1] YX_right[0] VDDP VSS INTCLKX_right / S013EELPSP_LEAFCELL_FPREDEC_YX
XI3 YA[0] YA[1] ACTRCLK ACTRCLKX YX[3] YX[2] YX[1] YX[0] VDDP VSS INTCLKX /  S013EELPSP_LEAFCELL_FPREDEC_YX
XI13 XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] XA[0] YA[1] YA[0] CEN CLK  S[1] S[0] VDDP VSS WEN / S013EELPSP_LEAFCELL_ESDA13
XI19 XA[3] XA[4] ACTRCLK_right ACTRCLKX_right PXA_right[3] PXA_right[2]  PXA_right[1] PXA_right[0] RDE VDDP VSS / S013EELPSP_LEAFCELL_PXA
XIPA XA[3] XA[4] ACTRCLK ACTRCLKX PXA[3] PXA[2] PXA[1] PXA[0] RDE VDDP VSS /  S013EELPSP_LEAFCELL_PXA
XI22 XA[7] XA[8] ACTRCLK_right ACTRCLKX_right PXC_right[3] PXC_right[2]  PXC_right[1] PXC_right[0] VDDP VSS / S013EELPSP_LEAFCELL_PX4
XI21 XA[5] XA[6] ACTRCLK_right ACTRCLKX_right PXB_right[3] PXB_right[2]  PXB_right[1] PXB_right[0] VDDP VSS / S013EELPSP_LEAFCELL_PX4
XI10 XA[5] XA[6] ACTRCLK ACTRCLKX PXB[3] PXB[2] PXB[1] PXB[0] VDDP VSS /  S013EELPSP_LEAFCELL_PX4
XI11 XA[7] XA[8] ACTRCLK ACTRCLKX PXC[3] PXC[2] PXC[1] PXC[0] VDDP VSS /  S013EELPSP_LEAFCELL_PX4
XI23 XA[0] XA[1] XA[2] ACTRCLK_right ACTRCLKX_right FCKX_right[7]  FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2]  FCKX_right[1] FCKX_right[0] VDDP VSS INTCLKX_right / S013EELPSP_LEAFCELL_FPREDEC
XIFPRE XA[0] XA[1] XA[2] ACTRCLK ACTRCLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4]  FCKX[3] FCKX[2] FCKX[1] FCKX[0] VDDP VSS INTCLKX / S013EELPSP_LEAFCELL_FPREDEC
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_YMUX8 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1]  BL[0] BLX[7] BLX[6] BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] DB DBX DIN  DINX VDDP VSS YS[7] YS[6] YS[5] YS[4] YS[3] YS[2] YS[1] YS[0]
*.PININFO DIN:I DINX:I YS[7]:I YS[6]:I YS[5]:I YS[4]:I YS[3]:I YS[2]:I YS[1]:I 
*.PININFO YS[0]:I BL[7]:B BL[6]:B BL[5]:B BL[4]:B BL[3]:B BL[2]:B BL[1]:B 
*.PININFO BL[0]:B BLX[7]:B BLX[6]:B BLX[5]:B BLX[4]:B BLX[3]:B BLX[2]:B 
*.PININFO BLX[1]:B BLX[0]:B DB:B DBX:B VDD:B VSS:B
XI11 BL[4] BLX[4] DB DBX DIN DINX VDDP VSS YS[4] / S013EELPSP_LEAFCELL_YMUXB
XI12 BL[5] BLX[5] DB DBX DIN DINX VDDP VSS YS[5] / S013EELPSP_LEAFCELL_YMUXB
XI13 BL[6] BLX[6] DB DBX DIN DINX VDDP VSS YS[6] / S013EELPSP_LEAFCELL_YMUXB
XI14 BL[7] BLX[7] DB DBX DIN DINX VDDP VSS YS[7] / S013EELPSP_LEAFCELL_YMUXB
XI3 BL[3] BLX[3] DB DBX DIN DINX VDDP VSS YS[3] / S013EELPSP_LEAFCELL_YMUXB
XI2 BL[2] BLX[2] DB DBX DIN DINX VDDP VSS YS[2] / S013EELPSP_LEAFCELL_YMUXB
XI1 BL[1] BLX[1] DB DBX DIN DINX VDDP VSS YS[1] / S013EELPSP_LEAFCELL_YMUXB
XI0 BL[0] BLX[0] DB DBX DIN DINX VDDP VSS YS[0] / S013EELPSP_LEAFCELL_YMUXB
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_YMX8SAWR_BW BL[7] BL[6] BL[5] BL[4] BL[3] BL[2]  BL[1] BL[0] BLX[7] BLX[6] BLX[5] BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] BWEN CLK  CLKX DATA DOUT SACK1 SACK4 VDDP VSS WE YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]  YX[1] YX[0]
*.PININFO BWEN:I CLK:I CLKX:I DATA:I SACK1:I SACK4:I WE:I YX[7]:I YX[6]:I 
*.PININFO YX[5]:I YX[4]:I YX[3]:I YX[2]:I YX[1]:I YX[0]:I DOUT:O BL[7]:B 
*.PININFO BL[6]:B BL[5]:B BL[4]:B BL[3]:B BL[2]:B BL[1]:B BL[0]:B BLX[7]:B 
*.PININFO BLX[6]:B BLX[5]:B BLX[4]:B BLX[3]:B BLX[2]:B BLX[1]:B BLX[0]:B VDD:B 
*.PININFO VSS:B
XIYMUX4 BL[7] BL[6] BL[5] BL[4] BL[3] BL[2] BL[1] BL[0] BLX[7] BLX[6] BLX[5]  BLX[4] BLX[3] BLX[2] BLX[1] BLX[0] DB DBX DIN DINX VDDP VSS net86[7] net86[6]  net86[5] net86[4] net86[3] net86[2] net86[1] net86[0] /  S013EELPSP_LEAFCELL_YMUX8
XISA DB DBX DOUT VDDP VSS SACK1 SACK4 / S013EELPSP_LEAFCELL_SA8
MN1 BWEN VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MN3 DATA VSS VSS VSS N15LL W=300.0n L=130.00n m=1
MP1 BWEN VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
MP3 DATA VDDP VDDP VDDP P15LL W=300.0n L=130.00n m=1
XI14[7] YX[7] VDDP VSS net86[7] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[6] YX[6] VDDP VSS net86[6] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[5] YX[5] VDDP VSS net86[5] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[4] YX[4] VDDP VSS net86[4] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[3] YX[3] VDDP VSS net86[3] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[2] YX[2] VDDP VSS net86[2] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[1] YX[1] VDDP VSS net86[1] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XI14[0] YX[0] VDDP VSS net86[0] / inv pl=130.00n pw=800.0n nl=130.00n nw=800.0n
XIDATAIN BWEN CLK CLKX DIN DATA DINX VDDP VSS WE / S013EELPSP_LEAFCELL_DATAIN
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_Logic_common_mode_Y8 ACTRCLK ACTRCLKX  ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX DCTRCLKX_right  DCTRCLK_right EMCLK FB_right FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2]  FCKX[1] FCKX[0] FCKX_right[7] FCKX_right[6] FCKX_right[5] FCKX_right[4]  FCKX_right[3] FCKX_right[2] FCKX_right[1] FCKX_right[0] INTCLKX  INTCLKX_right PXA[3] PXA[2] PXA[1] PXA[0] PXA_right[3] PXA_right[2]  PXA_right[1] PXA_right[0] PXB[3] PXB[2] PXB[1] PXB[0] PXB_right[3]  PXB_right[2] PXB_right[1] PXB_right[0] PXC[3] PXC[2] PXC[1] PXC[0]  PXC_right[3] PXC_right[2] PXC_right[1] PXC_right[0] RDE S[1] S[0] SACK1  SACK1_right SACK4 SACK4_right SM VDDP VMINE VSS WE WEN WE_right XA[8] XA[7]  XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] XA[0] YA[2] YA[1] YA[0] YX[7] YX[6]  YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] YX_right[7] YX_right[6] YX_right[5]  YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0]
*.PININFO CEN:I CLK:I FB_right:I RDE:I S[1]:I S[0]:I SM:I VMINE:I WEN:I 
*.PININFO XA[8]:I XA[7]:I XA[6]:I XA[5]:I XA[4]:I XA[3]:I XA[2]:I XA[1]:I 
*.PININFO XA[0]:I YA[2]:I YA[1]:I YA[0]:I ACTRCLK:O ACTRCLKX:O 
*.PININFO ACTRCLKX_right:O ACTRCLK_right:O DCTRCLK:O DCTRCLKX:O 
*.PININFO DCTRCLKX_right:O DCTRCLK_right:O EMCLK:O FCKX[7]:O FCKX[6]:O 
*.PININFO FCKX[5]:O FCKX[4]:O FCKX[3]:O FCKX[2]:O FCKX[1]:O FCKX[0]:O 
*.PININFO FCKX_right[7]:O FCKX_right[6]:O FCKX_right[5]:O FCKX_right[4]:O 
*.PININFO FCKX_right[3]:O FCKX_right[2]:O FCKX_right[1]:O FCKX_right[0]:O 
*.PININFO INTCLKX:O INTCLKX_right:O PXA[3]:O PXA[2]:O PXA[1]:O PXA[0]:O 
*.PININFO PXA_right[3]:O PXA_right[2]:O PXA_right[1]:O PXA_right[0]:O PXB[3]:O 
*.PININFO PXB[2]:O PXB[1]:O PXB[0]:O PXB_right[3]:O PXB_right[2]:O 
*.PININFO PXB_right[1]:O PXB_right[0]:O PXC[3]:O PXC[2]:O PXC[1]:O PXC[0]:O 
*.PININFO PXC_right[3]:O PXC_right[2]:O PXC_right[1]:O PXC_right[0]:O SACK1:O 
*.PININFO SACK1_right:O SACK4:O SACK4_right:O WE:O WE_right:O YX[7]:O YX[6]:O 
*.PININFO YX[5]:O YX[4]:O YX[3]:O YX[2]:O YX[1]:O YX[0]:O YX_right[7]:O 
*.PININFO YX_right[6]:O YX_right[5]:O YX_right[4]:O YX_right[3]:O 
*.PININFO YX_right[2]:O YX_right[1]:O YX_right[0]:O VDD:B VSS:B
XICLKDRV ACTRCLK ACTRCLKX ACTRCLKX_right ACTRCLK_right CEN CLK DCTRCLK DCTRCLKX  DCTRCLKX_right DCTRCLK_right EMCLK FB_right INTCLKX INTCLKX_right S[1] S[0]  SACK1 SACK1_right SACK4 SACK4_right SM VDDP VMINE VSS WE WEN WE_right /  S013EELPSP_LEAFCELL_CLKDRV_mode_V1
XI13 XA[8] XA[7] XA[6] XA[5] XA[4] XA[3] XA[2] XA[1] XA[0] YA[2] YA[1] YA[0] CEN CLK  S[1] S[0] VDDP VSS WEN / S013EELPSP_LEAFCELL_ESDA14
XI19 XA[3] XA[4] ACTRCLK_right ACTRCLKX_right PXA_right[3] PXA_right[2]  PXA_right[1] PXA_right[0] RDE VDDP VSS / S013EELPSP_LEAFCELL_PXA
XPA XA[3] XA[4] ACTRCLK ACTRCLKX PXA[3] PXA[2] PXA[1] PXA[0] RDE VDDP VSS /  S013EELPSP_LEAFCELL_PXA
XI22 XA[7] XA[8] ACTRCLK_right ACTRCLKX_right PXC_right[3] PXC_right[2]  PXC_right[1] PXC_right[0] VDDP VSS / S013EELPSP_LEAFCELL_PX4
XI21 XA[5] XA[6] ACTRCLK_right ACTRCLKX_right PXB_right[3] PXB_right[2]  PXB_right[1] PXB_right[0] VDDP VSS / S013EELPSP_LEAFCELL_PX4
XI10 XA[5] XA[6] ACTRCLK ACTRCLKX PXB[3] PXB[2] PXB[1] PXB[0] VDDP VSS /  S013EELPSP_LEAFCELL_PX4
XI11 XA[7] XA[8] ACTRCLK ACTRCLKX PXC[3] PXC[2] PXC[1] PXC[0] VDDP VSS /  S013EELPSP_LEAFCELL_PX4
XI26 YA[0] YA[1] YA[2] ACTRCLK_right ACTRCLKX_right YX_right[7] YX_right[6]  YX_right[5] YX_right[4] YX_right[3] YX_right[2] YX_right[1] YX_right[0] VDDP  VSS INTCLKX_right / S013EELPSP_LEAFCELL_FPREDEC
XI23 XA[0] XA[1] XA[2] ACTRCLK_right ACTRCLKX_right FCKX_right[7]  FCKX_right[6] FCKX_right[5] FCKX_right[4] FCKX_right[3] FCKX_right[2]  FCKX_right[1] FCKX_right[0] VDDP VSS INTCLKX_right / S013EELPSP_LEAFCELL_FPREDEC
XI25 YA[0] YA[1] YA[2] ACTRCLK ACTRCLKX YX[7] YX[6] YX[5] YX[4] YX[3] YX[2]  YX[1] YX[0] VDDP VSS INTCLKX / S013EELPSP_LEAFCELL_FPREDEC
XIFPRE XA[0] XA[1] XA[2] ACTRCLK ACTRCLKX FCKX[7] FCKX[6] FCKX[5] FCKX[4]  FCKX[3] FCKX[2] FCKX[1] FCKX[0] VDDP VSS INTCLKX / S013EELPSP_LEAFCELL_FPREDEC
.ENDS

.SUBCKT S013EELPSP_LEAFCELL_FDEC_right_V0P11 FCKX PABC PABCX VDDP VSS WLR
MM2 WLR net46 VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS net46 / inv pl=130.00n pw=2u nl=150.00n nw=1.5u
XI8 A VDDP VSS B / inv pl=130.00n pw=700.0n nl=130.00n nw=1u
XI114 A PABC PABCX VDDP VSS FCKX / tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
MM3 WLR net46 VDDP VDDP P15LL W=2.5u L=150.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_FDEC_left_V0P11 FCKX PABC PABCX VDDP VSS WLL
MM1 WLL C VSS VSS N15LL W=2u L=130.00n m=1
XI7 B VDDP VSS C / inv pl=130.00n pw=2u nl=150.00n nw=1.5u
XI8 A VDDP VSS B / inv pl=130.00n pw=700.0n nl=130.00n nw=1u
XI114 A PABC PABCX VDDP VSS FCKX / tgate pl=130.00n pw=800.0n nl=130.00n nw=1.2u
MM0 WLL C VDDP VDDP P15LL W=2.5u L=150.00n m=1
MP9 A PABC VDDP VDDP P15LL W=800.0n L=130.00n m=1
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_XDEC_right_V0P11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] 
+ FCKX[2] FCKX[1] FCKX[0] PXA PXB PXC VDDP VSS WLR[7] WLR[6] WLR[5] WLR[4] 
+ WLR[3] WLR[2] WLR[1] WLR[0]
*.PININFO FCKX[7]:I FCKX[6]:I FCKX[5]:I FCKX[4]:I FCKX[3]:I FCKX[2]:I 
*.PININFO FCKX[1]:I FCKX[0]:I PXA:I PXB:I PXC:I WLR[7]:O WLR[6]:O WLR[5]:O 
*.PININFO WLR[4]:O WLR[3]:O WLR[2]:O WLR[1]:O WLR[0]:O VDD:B VSS:B
XI156 PXA PXB PXC VDDP VSS net31 / nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLR[7] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLR[6] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLR[5] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLR[4] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLR[3] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLR[2] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLR[1] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLR[0] / S013EELPSP_LEAFCELL_FDEC_right_V0P11
XI111 net31 VDDP VSS PABC / inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS


.SUBCKT S013EELPSP_LEAFCELL_XDEC_left_V0P11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] 
+ FCKX[2] FCKX[1] FCKX[0] PXA PXB PXC VDDP VSS WLL[7] WLL[6] WLL[5] WLL[4] 
+ WLL[3] WLL[2] WLL[1] WLL[0]
*.PININFO FCKX[7]:I FCKX[6]:I FCKX[5]:I FCKX[4]:I FCKX[3]:I FCKX[2]:I 
*.PININFO FCKX[1]:I FCKX[0]:I PXA:I PXB:I PXC:I WLL[7]:O WLL[6]:O WLL[5]:O 
*.PININFO WLL[4]:O WLL[3]:O WLL[2]:O WLL[1]:O WLL[0]:O VDD:B VSS:B
XI156 PXA PXB PXC VDDP VSS net31 / nand3 pl=130.00n pw=1.0u nl=130.00n nw=2u
XFDEC[7] FCKX[7] PABC PABCX VDDP VSS WLL[7] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[6] FCKX[6] PABC PABCX VDDP VSS WLL[6] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[5] FCKX[5] PABC PABCX VDDP VSS WLL[5] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[4] FCKX[4] PABC PABCX VDDP VSS WLL[4] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[3] FCKX[3] PABC PABCX VDDP VSS WLL[3] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[2] FCKX[2] PABC PABCX VDDP VSS WLL[2] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[1] FCKX[1] PABC PABCX VDDP VSS WLL[1] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XFDEC[0] FCKX[0] PABC PABCX VDDP VSS WLL[0] / S013EELPSP_LEAFCELL_FDEC_left_V0P11
XI111 net31 VDDP VSS PABC / inv pl=130.00n pw=3u nl=130.00n nw=2u
XI112 PABC VDDP VSS PABCX / inv pl=130.00n pw=2u nl=130.00n nw=2u
.ENDS


